// This is the unpowered netlist.
module tiny_user_project (user_clock2,
    wb_clk_i,
    wb_rst_i,
    wbs_ack_o,
    wbs_cyc_i,
    wbs_stb_i,
    wbs_we_i,
    io_in,
    io_oeb,
    io_out,
    la_data_in,
    la_data_out,
    la_oenb,
    user_irq,
    wbs_adr_i,
    wbs_dat_i,
    wbs_dat_o,
    wbs_sel_i);
 input user_clock2;
 input wb_clk_i;
 input wb_rst_i;
 output wbs_ack_o;
 input wbs_cyc_i;
 input wbs_stb_i;
 input wbs_we_i;
 input [37:0] io_in;
 output [37:0] io_oeb;
 output [37:0] io_out;
 input [63:0] la_data_in;
 output [63:0] la_data_out;
 input [63:0] la_oenb;
 output [2:0] user_irq;
 input [31:0] wbs_adr_i;
 input [31:0] wbs_dat_i;
 output [31:0] wbs_dat_o;
 input [3:0] wbs_sel_i;

 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire net191;
 wire net190;
 wire net189;
 wire net188;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire net187;
 wire net186;
 wire net185;
 wire net184;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire net183;
 wire net182;
 wire net181;
 wire net180;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire _0656_;
 wire _0657_;
 wire _0658_;
 wire _0659_;
 wire _0660_;
 wire _0661_;
 wire _0662_;
 wire _0663_;
 wire _0664_;
 wire _0665_;
 wire _0666_;
 wire _0667_;
 wire _0668_;
 wire _0669_;
 wire _0670_;
 wire _0671_;
 wire _0672_;
 wire _0673_;
 wire _0674_;
 wire _0675_;
 wire _0676_;
 wire _0677_;
 wire _0678_;
 wire _0679_;
 wire _0680_;
 wire _0681_;
 wire _0682_;
 wire _0683_;
 wire _0684_;
 wire _0685_;
 wire _0686_;
 wire _0687_;
 wire _0688_;
 wire _0689_;
 wire _0690_;
 wire _0691_;
 wire _0692_;
 wire _0693_;
 wire _0694_;
 wire _0695_;
 wire _0696_;
 wire _0697_;
 wire _0698_;
 wire _0699_;
 wire _0700_;
 wire _0701_;
 wire _0702_;
 wire _0703_;
 wire _0704_;
 wire _0705_;
 wire _0706_;
 wire _0707_;
 wire _0708_;
 wire _0709_;
 wire _0710_;
 wire _0711_;
 wire _0712_;
 wire _0713_;
 wire _0714_;
 wire _0715_;
 wire _0716_;
 wire _0717_;
 wire _0718_;
 wire _0719_;
 wire _0720_;
 wire _0721_;
 wire _0722_;
 wire _0723_;
 wire _0724_;
 wire _0725_;
 wire _0726_;
 wire _0727_;
 wire _0728_;
 wire _0729_;
 wire _0730_;
 wire _0731_;
 wire _0732_;
 wire _0733_;
 wire _0734_;
 wire _0735_;
 wire _0736_;
 wire _0737_;
 wire _0738_;
 wire _0739_;
 wire _0740_;
 wire _0741_;
 wire _0742_;
 wire _0743_;
 wire _0744_;
 wire _0745_;
 wire _0746_;
 wire _0747_;
 wire _0748_;
 wire _0749_;
 wire _0750_;
 wire _0751_;
 wire _0752_;
 wire _0753_;
 wire _0754_;
 wire _0755_;
 wire _0756_;
 wire _0757_;
 wire _0758_;
 wire _0759_;
 wire _0760_;
 wire _0761_;
 wire _0762_;
 wire _0763_;
 wire _0764_;
 wire _0765_;
 wire _0766_;
 wire _0767_;
 wire _0768_;
 wire _0769_;
 wire _0770_;
 wire _0771_;
 wire _0772_;
 wire _0773_;
 wire _0774_;
 wire _0775_;
 wire _0776_;
 wire _0777_;
 wire _0778_;
 wire _0779_;
 wire _0780_;
 wire _0781_;
 wire _0782_;
 wire _0783_;
 wire _0784_;
 wire _0785_;
 wire _0786_;
 wire _0787_;
 wire _0788_;
 wire _0789_;
 wire _0790_;
 wire _0791_;
 wire _0792_;
 wire _0793_;
 wire _0794_;
 wire _0795_;
 wire _0796_;
 wire _0797_;
 wire _0798_;
 wire _0799_;
 wire _0800_;
 wire _0801_;
 wire _0802_;
 wire _0803_;
 wire _0804_;
 wire _0805_;
 wire _0806_;
 wire _0807_;
 wire _0808_;
 wire _0809_;
 wire _0810_;
 wire _0811_;
 wire _0812_;
 wire _0813_;
 wire _0814_;
 wire _0815_;
 wire _0816_;
 wire _0817_;
 wire _0818_;
 wire _0819_;
 wire _0820_;
 wire _0821_;
 wire _0822_;
 wire _0823_;
 wire _0824_;
 wire _0825_;
 wire _0826_;
 wire _0827_;
 wire _0828_;
 wire _0829_;
 wire _0830_;
 wire _0831_;
 wire _0832_;
 wire _0833_;
 wire _0834_;
 wire _0835_;
 wire _0836_;
 wire _0837_;
 wire _0838_;
 wire _0839_;
 wire _0840_;
 wire _0841_;
 wire _0842_;
 wire _0843_;
 wire _0844_;
 wire _0845_;
 wire _0846_;
 wire _0847_;
 wire _0848_;
 wire _0849_;
 wire _0850_;
 wire _0851_;
 wire _0852_;
 wire _0853_;
 wire _0854_;
 wire _0855_;
 wire _0856_;
 wire _0857_;
 wire _0858_;
 wire _0859_;
 wire _0860_;
 wire _0861_;
 wire _0862_;
 wire _0863_;
 wire _0864_;
 wire _0865_;
 wire _0866_;
 wire _0867_;
 wire _0868_;
 wire _0869_;
 wire _0870_;
 wire _0871_;
 wire _0872_;
 wire _0873_;
 wire _0874_;
 wire _0875_;
 wire _0876_;
 wire _0877_;
 wire _0878_;
 wire _0879_;
 wire _0880_;
 wire _0881_;
 wire _0882_;
 wire _0883_;
 wire _0884_;
 wire _0885_;
 wire _0886_;
 wire _0887_;
 wire _0888_;
 wire _0889_;
 wire _0890_;
 wire _0891_;
 wire _0892_;
 wire _0893_;
 wire _0894_;
 wire _0895_;
 wire _0896_;
 wire _0897_;
 wire _0898_;
 wire _0899_;
 wire _0900_;
 wire _0901_;
 wire _0902_;
 wire _0903_;
 wire _0904_;
 wire _0905_;
 wire _0906_;
 wire _0907_;
 wire _0908_;
 wire _0909_;
 wire _0910_;
 wire _0911_;
 wire _0912_;
 wire _0913_;
 wire _0914_;
 wire _0915_;
 wire _0916_;
 wire _0917_;
 wire _0918_;
 wire _0919_;
 wire _0920_;
 wire _0921_;
 wire _0922_;
 wire _0923_;
 wire _0924_;
 wire _0925_;
 wire _0926_;
 wire _0927_;
 wire _0928_;
 wire _0929_;
 wire _0930_;
 wire _0931_;
 wire _0932_;
 wire _0933_;
 wire _0934_;
 wire _0935_;
 wire _0936_;
 wire _0937_;
 wire _0938_;
 wire _0939_;
 wire _0940_;
 wire _0941_;
 wire _0942_;
 wire _0943_;
 wire _0944_;
 wire _0945_;
 wire _0946_;
 wire _0947_;
 wire _0948_;
 wire _0949_;
 wire _0950_;
 wire _0951_;
 wire _0952_;
 wire _0953_;
 wire _0954_;
 wire _0955_;
 wire _0956_;
 wire _0957_;
 wire _0958_;
 wire _0959_;
 wire _0960_;
 wire _0961_;
 wire _0962_;
 wire _0963_;
 wire _0964_;
 wire _0965_;
 wire _0966_;
 wire _0967_;
 wire _0968_;
 wire _0969_;
 wire _0970_;
 wire _0971_;
 wire _0972_;
 wire _0973_;
 wire _0974_;
 wire _0975_;
 wire _0976_;
 wire _0977_;
 wire _0978_;
 wire _0979_;
 wire _0980_;
 wire _0981_;
 wire _0982_;
 wire _0983_;
 wire _0984_;
 wire _0985_;
 wire _0986_;
 wire _0987_;
 wire _0988_;
 wire _0989_;
 wire _0990_;
 wire _0991_;
 wire _0992_;
 wire _0993_;
 wire _0994_;
 wire _0995_;
 wire _0996_;
 wire _0997_;
 wire _0998_;
 wire _0999_;
 wire _1000_;
 wire _1001_;
 wire _1002_;
 wire _1003_;
 wire _1004_;
 wire _1005_;
 wire _1006_;
 wire _1007_;
 wire _1008_;
 wire _1009_;
 wire _1010_;
 wire _1011_;
 wire _1012_;
 wire _1013_;
 wire _1014_;
 wire _1015_;
 wire _1016_;
 wire _1017_;
 wire _1018_;
 wire _1019_;
 wire _1020_;
 wire _1021_;
 wire _1022_;
 wire _1023_;
 wire _1024_;
 wire _1025_;
 wire _1026_;
 wire _1027_;
 wire _1028_;
 wire _1029_;
 wire _1030_;
 wire _1031_;
 wire _1032_;
 wire _1033_;
 wire _1034_;
 wire _1035_;
 wire _1036_;
 wire _1037_;
 wire _1038_;
 wire _1039_;
 wire _1040_;
 wire _1041_;
 wire _1042_;
 wire _1043_;
 wire _1044_;
 wire _1045_;
 wire _1046_;
 wire _1047_;
 wire _1048_;
 wire _1049_;
 wire _1050_;
 wire _1051_;
 wire _1052_;
 wire _1053_;
 wire _1054_;
 wire _1055_;
 wire _1056_;
 wire _1057_;
 wire _1058_;
 wire _1059_;
 wire _1060_;
 wire _1061_;
 wire _1062_;
 wire _1063_;
 wire _1064_;
 wire _1065_;
 wire _1066_;
 wire _1067_;
 wire _1068_;
 wire _1069_;
 wire _1070_;
 wire _1071_;
 wire _1072_;
 wire _1073_;
 wire _1074_;
 wire _1075_;
 wire _1076_;
 wire _1077_;
 wire _1078_;
 wire _1079_;
 wire _1080_;
 wire _1081_;
 wire _1082_;
 wire _1083_;
 wire _1084_;
 wire _1085_;
 wire _1086_;
 wire _1087_;
 wire _1088_;
 wire _1089_;
 wire _1090_;
 wire _1091_;
 wire _1092_;
 wire _1093_;
 wire _1094_;
 wire _1095_;
 wire _1096_;
 wire _1097_;
 wire _1098_;
 wire _1099_;
 wire _1100_;
 wire _1101_;
 wire _1102_;
 wire _1103_;
 wire _1104_;
 wire _1105_;
 wire _1106_;
 wire _1107_;
 wire _1108_;
 wire _1109_;
 wire _1110_;
 wire _1111_;
 wire _1112_;
 wire _1113_;
 wire _1114_;
 wire _1115_;
 wire _1116_;
 wire _1117_;
 wire _1118_;
 wire _1119_;
 wire _1120_;
 wire _1121_;
 wire _1122_;
 wire _1123_;
 wire _1124_;
 wire _1125_;
 wire _1126_;
 wire _1127_;
 wire _1128_;
 wire _1129_;
 wire _1130_;
 wire _1131_;
 wire _1132_;
 wire _1133_;
 wire _1134_;
 wire _1135_;
 wire _1136_;
 wire _1137_;
 wire _1138_;
 wire _1139_;
 wire _1140_;
 wire _1141_;
 wire _1142_;
 wire _1143_;
 wire _1144_;
 wire _1145_;
 wire _1146_;
 wire _1147_;
 wire _1148_;
 wire _1149_;
 wire _1150_;
 wire _1151_;
 wire _1152_;
 wire _1153_;
 wire _1154_;
 wire _1155_;
 wire _1156_;
 wire _1157_;
 wire _1158_;
 wire _1159_;
 wire _1160_;
 wire _1161_;
 wire _1162_;
 wire _1163_;
 wire _1164_;
 wire _1165_;
 wire _1166_;
 wire _1167_;
 wire _1168_;
 wire _1169_;
 wire _1170_;
 wire _1171_;
 wire _1172_;
 wire _1173_;
 wire _1174_;
 wire _1175_;
 wire _1176_;
 wire _1177_;
 wire _1178_;
 wire _1179_;
 wire _1180_;
 wire _1181_;
 wire _1182_;
 wire _1183_;
 wire _1184_;
 wire _1185_;
 wire _1186_;
 wire _1187_;
 wire _1188_;
 wire _1189_;
 wire _1190_;
 wire _1191_;
 wire _1192_;
 wire _1193_;
 wire _1194_;
 wire _1195_;
 wire _1196_;
 wire _1197_;
 wire _1198_;
 wire _1199_;
 wire _1200_;
 wire _1201_;
 wire _1202_;
 wire _1203_;
 wire _1204_;
 wire _1205_;
 wire _1206_;
 wire _1207_;
 wire _1208_;
 wire _1209_;
 wire _1210_;
 wire _1211_;
 wire _1212_;
 wire _1213_;
 wire _1214_;
 wire _1215_;
 wire _1216_;
 wire _1217_;
 wire _1218_;
 wire _1219_;
 wire _1220_;
 wire _1221_;
 wire _1222_;
 wire _1223_;
 wire _1224_;
 wire _1225_;
 wire _1226_;
 wire _1227_;
 wire _1228_;
 wire _1229_;
 wire _1230_;
 wire _1231_;
 wire _1232_;
 wire _1233_;
 wire _1234_;
 wire _1235_;
 wire _1236_;
 wire _1237_;
 wire _1238_;
 wire _1239_;
 wire _1240_;
 wire _1241_;
 wire _1242_;
 wire _1243_;
 wire _1244_;
 wire _1245_;
 wire _1246_;
 wire _1247_;
 wire _1248_;
 wire _1249_;
 wire _1250_;
 wire _1251_;
 wire _1252_;
 wire _1253_;
 wire _1254_;
 wire _1255_;
 wire _1256_;
 wire _1257_;
 wire _1258_;
 wire _1259_;
 wire _1260_;
 wire _1261_;
 wire _1262_;
 wire _1263_;
 wire _1264_;
 wire _1265_;
 wire _1266_;
 wire _1267_;
 wire _1268_;
 wire _1269_;
 wire _1270_;
 wire _1271_;
 wire _1272_;
 wire _1273_;
 wire _1274_;
 wire _1275_;
 wire _1276_;
 wire _1277_;
 wire _1278_;
 wire _1279_;
 wire _1280_;
 wire _1281_;
 wire _1282_;
 wire _1283_;
 wire _1284_;
 wire _1285_;
 wire _1286_;
 wire _1287_;
 wire _1288_;
 wire _1289_;
 wire _1290_;
 wire _1291_;
 wire _1292_;
 wire _1293_;
 wire _1294_;
 wire _1295_;
 wire _1296_;
 wire _1297_;
 wire _1298_;
 wire _1299_;
 wire _1300_;
 wire _1301_;
 wire _1302_;
 wire _1303_;
 wire _1304_;
 wire _1305_;
 wire _1306_;
 wire _1307_;
 wire _1308_;
 wire _1309_;
 wire _1310_;
 wire _1311_;
 wire _1312_;
 wire _1313_;
 wire _1314_;
 wire _1315_;
 wire _1316_;
 wire _1317_;
 wire _1318_;
 wire _1319_;
 wire _1320_;
 wire _1321_;
 wire _1322_;
 wire _1323_;
 wire _1324_;
 wire _1325_;
 wire _1326_;
 wire _1327_;
 wire _1328_;
 wire _1329_;
 wire _1330_;
 wire _1331_;
 wire _1332_;
 wire _1333_;
 wire _1334_;
 wire _1335_;
 wire _1336_;
 wire _1337_;
 wire _1338_;
 wire _1339_;
 wire _1340_;
 wire _1341_;
 wire _1342_;
 wire _1343_;
 wire _1344_;
 wire _1345_;
 wire _1346_;
 wire _1347_;
 wire _1348_;
 wire _1349_;
 wire _1350_;
 wire _1351_;
 wire _1352_;
 wire _1353_;
 wire _1354_;
 wire _1355_;
 wire _1356_;
 wire _1357_;
 wire _1358_;
 wire _1359_;
 wire _1360_;
 wire _1361_;
 wire _1362_;
 wire _1363_;
 wire _1364_;
 wire _1365_;
 wire _1366_;
 wire _1367_;
 wire _1368_;
 wire _1369_;
 wire _1370_;
 wire _1371_;
 wire _1372_;
 wire _1373_;
 wire _1374_;
 wire _1375_;
 wire _1376_;
 wire _1377_;
 wire _1378_;
 wire _1379_;
 wire _1380_;
 wire _1381_;
 wire _1382_;
 wire _1383_;
 wire _1384_;
 wire _1385_;
 wire _1386_;
 wire _1387_;
 wire _1388_;
 wire _1389_;
 wire _1390_;
 wire _1391_;
 wire _1392_;
 wire _1393_;
 wire _1394_;
 wire _1395_;
 wire _1396_;
 wire _1397_;
 wire _1398_;
 wire _1399_;
 wire _1400_;
 wire _1401_;
 wire _1402_;
 wire _1403_;
 wire _1404_;
 wire _1405_;
 wire _1406_;
 wire _1407_;
 wire _1408_;
 wire _1409_;
 wire _1410_;
 wire _1411_;
 wire _1412_;
 wire _1413_;
 wire _1414_;
 wire _1415_;
 wire _1416_;
 wire _1417_;
 wire _1418_;
 wire _1419_;
 wire _1420_;
 wire _1421_;
 wire _1422_;
 wire _1423_;
 wire _1424_;
 wire _1425_;
 wire _1426_;
 wire _1427_;
 wire _1428_;
 wire _1429_;
 wire _1430_;
 wire _1431_;
 wire _1432_;
 wire _1433_;
 wire _1434_;
 wire _1435_;
 wire _1436_;
 wire _1437_;
 wire _1438_;
 wire _1439_;
 wire _1440_;
 wire _1441_;
 wire _1442_;
 wire _1443_;
 wire _1444_;
 wire _1445_;
 wire _1446_;
 wire _1447_;
 wire _1448_;
 wire _1449_;
 wire _1450_;
 wire _1451_;
 wire _1452_;
 wire _1453_;
 wire _1454_;
 wire _1455_;
 wire _1456_;
 wire _1457_;
 wire _1458_;
 wire _1459_;
 wire _1460_;
 wire _1461_;
 wire _1462_;
 wire _1463_;
 wire _1464_;
 wire _1465_;
 wire _1466_;
 wire _1467_;
 wire _1468_;
 wire _1469_;
 wire _1470_;
 wire _1471_;
 wire _1472_;
 wire _1473_;
 wire _1474_;
 wire _1475_;
 wire _1476_;
 wire _1477_;
 wire _1478_;
 wire _1479_;
 wire _1480_;
 wire _1481_;
 wire _1482_;
 wire _1483_;
 wire _1484_;
 wire _1485_;
 wire _1486_;
 wire _1487_;
 wire _1488_;
 wire _1489_;
 wire _1490_;
 wire _1491_;
 wire _1492_;
 wire _1493_;
 wire _1494_;
 wire _1495_;
 wire _1496_;
 wire _1497_;
 wire _1498_;
 wire _1499_;
 wire _1500_;
 wire _1501_;
 wire _1502_;
 wire _1503_;
 wire _1504_;
 wire _1505_;
 wire _1506_;
 wire _1507_;
 wire _1508_;
 wire _1509_;
 wire _1510_;
 wire _1511_;
 wire _1512_;
 wire _1513_;
 wire _1514_;
 wire _1515_;
 wire _1516_;
 wire _1517_;
 wire _1518_;
 wire _1519_;
 wire _1520_;
 wire _1521_;
 wire _1522_;
 wire _1523_;
 wire _1524_;
 wire _1525_;
 wire _1526_;
 wire _1527_;
 wire _1528_;
 wire _1529_;
 wire _1530_;
 wire _1531_;
 wire _1532_;
 wire _1533_;
 wire _1534_;
 wire _1535_;
 wire _1536_;
 wire _1537_;
 wire _1538_;
 wire _1539_;
 wire _1540_;
 wire _1541_;
 wire _1542_;
 wire _1543_;
 wire _1544_;
 wire _1545_;
 wire _1546_;
 wire _1547_;
 wire _1548_;
 wire _1549_;
 wire _1550_;
 wire _1551_;
 wire _1552_;
 wire _1553_;
 wire _1554_;
 wire _1555_;
 wire _1556_;
 wire _1557_;
 wire _1558_;
 wire _1559_;
 wire _1560_;
 wire _1561_;
 wire _1562_;
 wire _1563_;
 wire _1564_;
 wire _1565_;
 wire _1566_;
 wire _1567_;
 wire _1568_;
 wire _1569_;
 wire _1570_;
 wire _1571_;
 wire _1572_;
 wire _1573_;
 wire _1574_;
 wire _1575_;
 wire _1576_;
 wire _1577_;
 wire _1578_;
 wire _1579_;
 wire _1580_;
 wire _1581_;
 wire _1582_;
 wire _1583_;
 wire _1584_;
 wire _1585_;
 wire _1586_;
 wire _1587_;
 wire _1588_;
 wire _1589_;
 wire _1590_;
 wire _1591_;
 wire _1592_;
 wire _1593_;
 wire _1594_;
 wire _1595_;
 wire _1596_;
 wire _1597_;
 wire _1598_;
 wire _1599_;
 wire _1600_;
 wire _1601_;
 wire _1602_;
 wire _1603_;
 wire _1604_;
 wire _1605_;
 wire _1606_;
 wire _1607_;
 wire _1608_;
 wire _1609_;
 wire _1610_;
 wire _1611_;
 wire _1612_;
 wire _1613_;
 wire _1614_;
 wire _1615_;
 wire _1616_;
 wire _1617_;
 wire _1618_;
 wire _1619_;
 wire _1620_;
 wire _1621_;
 wire _1622_;
 wire _1623_;
 wire _1624_;
 wire _1625_;
 wire _1626_;
 wire _1627_;
 wire _1628_;
 wire _1629_;
 wire _1630_;
 wire _1631_;
 wire _1632_;
 wire _1633_;
 wire _1634_;
 wire _1635_;
 wire _1636_;
 wire _1637_;
 wire _1638_;
 wire _1639_;
 wire _1640_;
 wire _1641_;
 wire _1642_;
 wire _1643_;
 wire _1644_;
 wire _1645_;
 wire _1646_;
 wire _1647_;
 wire _1648_;
 wire _1649_;
 wire _1650_;
 wire _1651_;
 wire _1652_;
 wire _1653_;
 wire _1654_;
 wire _1655_;
 wire _1656_;
 wire _1657_;
 wire _1658_;
 wire _1659_;
 wire _1660_;
 wire _1661_;
 wire _1662_;
 wire _1663_;
 wire _1664_;
 wire _1665_;
 wire _1666_;
 wire _1667_;
 wire _1668_;
 wire _1669_;
 wire _1670_;
 wire _1671_;
 wire _1672_;
 wire _1673_;
 wire _1674_;
 wire _1675_;
 wire _1676_;
 wire _1677_;
 wire _1678_;
 wire _1679_;
 wire _1680_;
 wire _1681_;
 wire _1682_;
 wire _1683_;
 wire _1684_;
 wire _1685_;
 wire _1686_;
 wire _1687_;
 wire _1688_;
 wire _1689_;
 wire _1690_;
 wire _1691_;
 wire _1692_;
 wire _1693_;
 wire _1694_;
 wire _1695_;
 wire _1696_;
 wire _1697_;
 wire _1698_;
 wire _1699_;
 wire _1700_;
 wire _1701_;
 wire _1702_;
 wire _1703_;
 wire _1704_;
 wire _1705_;
 wire _1706_;
 wire _1707_;
 wire _1708_;
 wire _1709_;
 wire _1710_;
 wire _1711_;
 wire _1712_;
 wire _1713_;
 wire _1714_;
 wire _1715_;
 wire _1716_;
 wire _1717_;
 wire _1718_;
 wire _1719_;
 wire _1720_;
 wire _1721_;
 wire _1722_;
 wire _1723_;
 wire _1724_;
 wire _1725_;
 wire _1726_;
 wire _1727_;
 wire _1728_;
 wire _1729_;
 wire _1730_;
 wire _1731_;
 wire _1732_;
 wire _1733_;
 wire _1734_;
 wire _1735_;
 wire _1736_;
 wire _1737_;
 wire _1738_;
 wire _1739_;
 wire _1740_;
 wire _1741_;
 wire _1742_;
 wire _1743_;
 wire _1744_;
 wire _1745_;
 wire _1746_;
 wire _1747_;
 wire _1748_;
 wire _1749_;
 wire _1750_;
 wire _1751_;
 wire _1752_;
 wire _1753_;
 wire _1754_;
 wire _1755_;
 wire _1756_;
 wire _1757_;
 wire _1758_;
 wire _1759_;
 wire _1760_;
 wire _1761_;
 wire _1762_;
 wire _1763_;
 wire _1764_;
 wire _1765_;
 wire _1766_;
 wire _1767_;
 wire _1768_;
 wire _1769_;
 wire _1770_;
 wire _1771_;
 wire _1772_;
 wire _1773_;
 wire _1774_;
 wire _1775_;
 wire _1776_;
 wire _1777_;
 wire _1778_;
 wire _1779_;
 wire _1780_;
 wire _1781_;
 wire _1782_;
 wire _1783_;
 wire _1784_;
 wire _1785_;
 wire _1786_;
 wire _1787_;
 wire _1788_;
 wire _1789_;
 wire _1790_;
 wire _1791_;
 wire _1792_;
 wire _1793_;
 wire _1794_;
 wire _1795_;
 wire _1796_;
 wire _1797_;
 wire _1798_;
 wire _1799_;
 wire _1800_;
 wire _1801_;
 wire _1802_;
 wire _1803_;
 wire _1804_;
 wire _1805_;
 wire _1806_;
 wire _1807_;
 wire _1808_;
 wire _1809_;
 wire _1810_;
 wire _1811_;
 wire _1812_;
 wire _1813_;
 wire _1814_;
 wire _1815_;
 wire _1816_;
 wire _1817_;
 wire _1818_;
 wire _1819_;
 wire _1820_;
 wire _1821_;
 wire _1822_;
 wire _1823_;
 wire _1824_;
 wire _1825_;
 wire _1826_;
 wire _1827_;
 wire _1828_;
 wire _1829_;
 wire _1830_;
 wire _1831_;
 wire _1832_;
 wire _1833_;
 wire _1834_;
 wire _1835_;
 wire _1836_;
 wire _1837_;
 wire _1838_;
 wire _1839_;
 wire _1840_;
 wire _1841_;
 wire _1842_;
 wire _1843_;
 wire _1844_;
 wire _1845_;
 wire _1846_;
 wire _1847_;
 wire _1848_;
 wire _1849_;
 wire _1850_;
 wire _1851_;
 wire _1852_;
 wire _1853_;
 wire _1854_;
 wire _1855_;
 wire _1856_;
 wire _1857_;
 wire _1858_;
 wire _1859_;
 wire _1860_;
 wire _1861_;
 wire _1862_;
 wire _1863_;
 wire _1864_;
 wire _1865_;
 wire _1866_;
 wire _1867_;
 wire _1868_;
 wire _1869_;
 wire _1870_;
 wire _1871_;
 wire _1872_;
 wire _1873_;
 wire _1874_;
 wire _1875_;
 wire _1876_;
 wire _1877_;
 wire _1878_;
 wire _1879_;
 wire _1880_;
 wire _1881_;
 wire _1882_;
 wire _1883_;
 wire _1884_;
 wire _1885_;
 wire _1886_;
 wire _1887_;
 wire _1888_;
 wire _1889_;
 wire _1890_;
 wire _1891_;
 wire _1892_;
 wire _1893_;
 wire _1894_;
 wire _1895_;
 wire _1896_;
 wire _1897_;
 wire _1898_;
 wire _1899_;
 wire _1900_;
 wire _1901_;
 wire _1902_;
 wire _1903_;
 wire _1904_;
 wire _1905_;
 wire _1906_;
 wire _1907_;
 wire _1908_;
 wire _1909_;
 wire _1910_;
 wire _1911_;
 wire _1912_;
 wire _1913_;
 wire _1914_;
 wire _1915_;
 wire _1916_;
 wire _1917_;
 wire _1918_;
 wire _1919_;
 wire _1920_;
 wire _1921_;
 wire _1922_;
 wire _1923_;
 wire _1924_;
 wire _1925_;
 wire _1926_;
 wire _1927_;
 wire _1928_;
 wire _1929_;
 wire _1930_;
 wire _1931_;
 wire _1932_;
 wire _1933_;
 wire _1934_;
 wire _1935_;
 wire _1936_;
 wire _1937_;
 wire _1938_;
 wire _1939_;
 wire _1940_;
 wire _1941_;
 wire _1942_;
 wire _1943_;
 wire _1944_;
 wire _1945_;
 wire _1946_;
 wire _1947_;
 wire _1948_;
 wire _1949_;
 wire _1950_;
 wire _1951_;
 wire _1952_;
 wire _1953_;
 wire _1954_;
 wire _1955_;
 wire _1956_;
 wire _1957_;
 wire _1958_;
 wire _1959_;
 wire _1960_;
 wire _1961_;
 wire _1962_;
 wire _1963_;
 wire _1964_;
 wire _1965_;
 wire _1966_;
 wire _1967_;
 wire _1968_;
 wire _1969_;
 wire _1970_;
 wire _1971_;
 wire _1972_;
 wire _1973_;
 wire _1974_;
 wire _1975_;
 wire _1976_;
 wire _1977_;
 wire _1978_;
 wire _1979_;
 wire _1980_;
 wire _1981_;
 wire _1982_;
 wire _1983_;
 wire _1984_;
 wire _1985_;
 wire _1986_;
 wire _1987_;
 wire _1988_;
 wire _1989_;
 wire _1990_;
 wire _1991_;
 wire _1992_;
 wire _1993_;
 wire _1994_;
 wire _1995_;
 wire _1996_;
 wire _1997_;
 wire _1998_;
 wire _1999_;
 wire _2000_;
 wire _2001_;
 wire _2002_;
 wire _2003_;
 wire _2004_;
 wire _2005_;
 wire _2006_;
 wire _2007_;
 wire _2008_;
 wire _2009_;
 wire _2010_;
 wire _2011_;
 wire _2012_;
 wire _2013_;
 wire _2014_;
 wire _2015_;
 wire _2016_;
 wire _2017_;
 wire _2018_;
 wire _2019_;
 wire _2020_;
 wire _2021_;
 wire _2022_;
 wire _2023_;
 wire _2024_;
 wire _2025_;
 wire _2026_;
 wire _2027_;
 wire _2028_;
 wire _2029_;
 wire _2030_;
 wire _2031_;
 wire _2032_;
 wire _2033_;
 wire _2034_;
 wire _2035_;
 wire _2036_;
 wire _2037_;
 wire _2038_;
 wire _2039_;
 wire _2040_;
 wire _2041_;
 wire _2042_;
 wire _2043_;
 wire _2044_;
 wire _2045_;
 wire _2046_;
 wire _2047_;
 wire _2048_;
 wire _2049_;
 wire _2050_;
 wire _2051_;
 wire _2052_;
 wire _2053_;
 wire _2054_;
 wire _2055_;
 wire _2056_;
 wire _2057_;
 wire _2058_;
 wire _2059_;
 wire _2060_;
 wire _2061_;
 wire _2062_;
 wire _2063_;
 wire _2064_;
 wire _2065_;
 wire _2066_;
 wire _2067_;
 wire _2068_;
 wire _2069_;
 wire _2070_;
 wire _2071_;
 wire _2072_;
 wire _2073_;
 wire _2074_;
 wire _2075_;
 wire _2076_;
 wire _2077_;
 wire _2078_;
 wire _2079_;
 wire _2080_;
 wire _2081_;
 wire _2082_;
 wire _2083_;
 wire _2084_;
 wire _2085_;
 wire _2086_;
 wire _2087_;
 wire _2088_;
 wire _2089_;
 wire _2090_;
 wire _2091_;
 wire _2092_;
 wire _2093_;
 wire _2094_;
 wire _2095_;
 wire _2096_;
 wire _2097_;
 wire _2098_;
 wire _2099_;
 wire _2100_;
 wire _2101_;
 wire _2102_;
 wire _2103_;
 wire _2104_;
 wire _2105_;
 wire _2106_;
 wire _2107_;
 wire _2108_;
 wire _2109_;
 wire _2110_;
 wire _2111_;
 wire _2112_;
 wire _2113_;
 wire _2114_;
 wire _2115_;
 wire _2116_;
 wire _2117_;
 wire _2118_;
 wire _2119_;
 wire _2120_;
 wire _2121_;
 wire _2122_;
 wire _2123_;
 wire _2124_;
 wire _2125_;
 wire _2126_;
 wire _2127_;
 wire _2128_;
 wire _2129_;
 wire _2130_;
 wire _2131_;
 wire _2132_;
 wire _2133_;
 wire _2134_;
 wire _2135_;
 wire _2136_;
 wire _2137_;
 wire _2138_;
 wire _2139_;
 wire _2140_;
 wire _2141_;
 wire _2142_;
 wire _2143_;
 wire _2144_;
 wire _2145_;
 wire _2146_;
 wire _2147_;
 wire _2148_;
 wire _2149_;
 wire _2150_;
 wire _2151_;
 wire _2152_;
 wire _2153_;
 wire _2154_;
 wire _2155_;
 wire _2156_;
 wire _2157_;
 wire _2158_;
 wire _2159_;
 wire _2160_;
 wire _2161_;
 wire _2162_;
 wire _2163_;
 wire _2164_;
 wire _2165_;
 wire _2166_;
 wire _2167_;
 wire _2168_;
 wire _2169_;
 wire _2170_;
 wire _2171_;
 wire _2172_;
 wire _2173_;
 wire _2174_;
 wire _2175_;
 wire _2176_;
 wire _2177_;
 wire _2178_;
 wire _2179_;
 wire _2180_;
 wire _2181_;
 wire _2182_;
 wire _2183_;
 wire _2184_;
 wire _2185_;
 wire _2186_;
 wire _2187_;
 wire _2188_;
 wire _2189_;
 wire _2190_;
 wire _2191_;
 wire _2192_;
 wire _2193_;
 wire _2194_;
 wire _2195_;
 wire _2196_;
 wire _2197_;
 wire _2198_;
 wire _2199_;
 wire _2200_;
 wire _2201_;
 wire _2202_;
 wire _2203_;
 wire _2204_;
 wire _2205_;
 wire _2206_;
 wire _2207_;
 wire _2208_;
 wire _2209_;
 wire _2210_;
 wire _2211_;
 wire _2212_;
 wire _2213_;
 wire _2214_;
 wire _2215_;
 wire _2216_;
 wire _2217_;
 wire _2218_;
 wire _2219_;
 wire _2220_;
 wire _2221_;
 wire _2222_;
 wire _2223_;
 wire _2224_;
 wire _2225_;
 wire _2226_;
 wire _2227_;
 wire _2228_;
 wire _2229_;
 wire _2230_;
 wire _2231_;
 wire _2232_;
 wire _2233_;
 wire _2234_;
 wire _2235_;
 wire _2236_;
 wire _2237_;
 wire _2238_;
 wire _2239_;
 wire _2240_;
 wire _2241_;
 wire _2242_;
 wire _2243_;
 wire _2244_;
 wire _2245_;
 wire _2246_;
 wire _2247_;
 wire _2248_;
 wire _2249_;
 wire _2250_;
 wire _2251_;
 wire _2252_;
 wire _2253_;
 wire _2254_;
 wire _2255_;
 wire _2256_;
 wire _2257_;
 wire _2258_;
 wire _2259_;
 wire _2260_;
 wire _2261_;
 wire _2262_;
 wire _2263_;
 wire _2264_;
 wire _2265_;
 wire _2266_;
 wire _2267_;
 wire _2268_;
 wire _2269_;
 wire _2270_;
 wire _2271_;
 wire _2272_;
 wire _2273_;
 wire _2274_;
 wire _2275_;
 wire _2276_;
 wire _2277_;
 wire _2278_;
 wire _2279_;
 wire _2280_;
 wire _2281_;
 wire _2282_;
 wire _2283_;
 wire _2284_;
 wire _2285_;
 wire _2286_;
 wire _2287_;
 wire _2288_;
 wire _2289_;
 wire _2290_;
 wire _2291_;
 wire _2292_;
 wire _2293_;
 wire _2294_;
 wire _2295_;
 wire _2296_;
 wire _2297_;
 wire _2298_;
 wire _2299_;
 wire _2300_;
 wire _2301_;
 wire _2302_;
 wire _2303_;
 wire _2304_;
 wire _2305_;
 wire _2306_;
 wire _2307_;
 wire _2308_;
 wire _2309_;
 wire _2310_;
 wire _2311_;
 wire _2312_;
 wire _2313_;
 wire _2314_;
 wire _2315_;
 wire _2316_;
 wire _2317_;
 wire _2318_;
 wire _2319_;
 wire _2320_;
 wire _2321_;
 wire _2322_;
 wire _2323_;
 wire _2324_;
 wire _2325_;
 wire _2326_;
 wire _2327_;
 wire _2328_;
 wire _2329_;
 wire _2330_;
 wire _2331_;
 wire _2332_;
 wire _2333_;
 wire _2334_;
 wire _2335_;
 wire _2336_;
 wire _2337_;
 wire _2338_;
 wire _2339_;
 wire _2340_;
 wire _2341_;
 wire _2342_;
 wire _2343_;
 wire _2344_;
 wire _2345_;
 wire _2346_;
 wire _2347_;
 wire _2348_;
 wire _2349_;
 wire _2350_;
 wire _2351_;
 wire _2352_;
 wire _2353_;
 wire _2354_;
 wire _2355_;
 wire _2356_;
 wire _2357_;
 wire _2358_;
 wire _2359_;
 wire _2360_;
 wire _2361_;
 wire _2362_;
 wire _2363_;
 wire _2364_;
 wire _2365_;
 wire _2366_;
 wire _2367_;
 wire _2368_;
 wire _2369_;
 wire _2370_;
 wire _2371_;
 wire _2372_;
 wire _2373_;
 wire _2374_;
 wire _2375_;
 wire _2376_;
 wire _2377_;
 wire _2378_;
 wire _2379_;
 wire _2380_;
 wire _2381_;
 wire _2382_;
 wire _2383_;
 wire _2384_;
 wire _2385_;
 wire _2386_;
 wire _2387_;
 wire _2388_;
 wire _2389_;
 wire _2390_;
 wire _2391_;
 wire _2392_;
 wire _2393_;
 wire _2394_;
 wire _2395_;
 wire _2396_;
 wire _2397_;
 wire _2398_;
 wire _2399_;
 wire _2400_;
 wire _2401_;
 wire _2402_;
 wire _2403_;
 wire _2404_;
 wire _2405_;
 wire _2406_;
 wire _2407_;
 wire _2408_;
 wire _2409_;
 wire _2410_;
 wire _2411_;
 wire _2412_;
 wire _2413_;
 wire _2414_;
 wire _2415_;
 wire _2416_;
 wire _2417_;
 wire _2418_;
 wire _2419_;
 wire _2420_;
 wire _2421_;
 wire _2422_;
 wire _2423_;
 wire _2424_;
 wire _2425_;
 wire _2426_;
 wire _2427_;
 wire _2428_;
 wire _2429_;
 wire _2430_;
 wire _2431_;
 wire _2432_;
 wire _2433_;
 wire _2434_;
 wire _2435_;
 wire _2436_;
 wire _2437_;
 wire _2438_;
 wire _2439_;
 wire _2440_;
 wire _2441_;
 wire _2442_;
 wire _2443_;
 wire _2444_;
 wire _2445_;
 wire _2446_;
 wire _2447_;
 wire _2448_;
 wire _2449_;
 wire _2450_;
 wire _2451_;
 wire _2452_;
 wire _2453_;
 wire _2454_;
 wire _2455_;
 wire _2456_;
 wire _2457_;
 wire _2458_;
 wire _2459_;
 wire _2460_;
 wire _2461_;
 wire _2462_;
 wire _2463_;
 wire _2464_;
 wire _2465_;
 wire _2466_;
 wire _2467_;
 wire _2468_;
 wire _2469_;
 wire _2470_;
 wire _2471_;
 wire _2472_;
 wire _2473_;
 wire _2474_;
 wire _2475_;
 wire _2476_;
 wire _2477_;
 wire _2478_;
 wire _2479_;
 wire _2480_;
 wire _2481_;
 wire _2482_;
 wire _2483_;
 wire _2484_;
 wire _2485_;
 wire _2486_;
 wire _2487_;
 wire _2488_;
 wire _2489_;
 wire _2490_;
 wire _2491_;
 wire _2492_;
 wire _2493_;
 wire _2494_;
 wire _2495_;
 wire _2496_;
 wire _2497_;
 wire _2498_;
 wire _2499_;
 wire _2500_;
 wire _2501_;
 wire _2502_;
 wire _2503_;
 wire _2504_;
 wire _2505_;
 wire _2506_;
 wire _2507_;
 wire _2508_;
 wire _2509_;
 wire _2510_;
 wire _2511_;
 wire _2512_;
 wire _2513_;
 wire _2514_;
 wire _2515_;
 wire _2516_;
 wire _2517_;
 wire _2518_;
 wire _2519_;
 wire _2520_;
 wire _2521_;
 wire _2522_;
 wire _2523_;
 wire _2524_;
 wire _2525_;
 wire _2526_;
 wire _2527_;
 wire _2528_;
 wire _2529_;
 wire _2530_;
 wire _2531_;
 wire _2532_;
 wire _2533_;
 wire _2534_;
 wire _2535_;
 wire _2536_;
 wire _2537_;
 wire _2538_;
 wire _2539_;
 wire _2540_;
 wire _2541_;
 wire _2542_;
 wire _2543_;
 wire _2544_;
 wire _2545_;
 wire _2546_;
 wire _2547_;
 wire _2548_;
 wire _2549_;
 wire _2550_;
 wire _2551_;
 wire _2552_;
 wire _2553_;
 wire _2554_;
 wire _2555_;
 wire _2556_;
 wire _2557_;
 wire _2558_;
 wire _2559_;
 wire _2560_;
 wire _2561_;
 wire _2562_;
 wire _2563_;
 wire _2564_;
 wire _2565_;
 wire _2566_;
 wire _2567_;
 wire _2568_;
 wire _2569_;
 wire _2570_;
 wire _2571_;
 wire _2572_;
 wire _2573_;
 wire _2574_;
 wire _2575_;
 wire _2576_;
 wire _2577_;
 wire _2578_;
 wire _2579_;
 wire _2580_;
 wire _2581_;
 wire _2582_;
 wire _2583_;
 wire _2584_;
 wire _2585_;
 wire _2586_;
 wire _2587_;
 wire _2588_;
 wire _2589_;
 wire _2590_;
 wire _2591_;
 wire _2592_;
 wire _2593_;
 wire _2594_;
 wire _2595_;
 wire _2596_;
 wire _2597_;
 wire _2598_;
 wire _2599_;
 wire _2600_;
 wire _2601_;
 wire _2602_;
 wire _2603_;
 wire _2604_;
 wire _2605_;
 wire _2606_;
 wire _2607_;
 wire _2608_;
 wire _2609_;
 wire _2610_;
 wire _2611_;
 wire _2612_;
 wire _2613_;
 wire _2614_;
 wire _2615_;
 wire _2616_;
 wire _2617_;
 wire _2618_;
 wire _2619_;
 wire _2620_;
 wire _2621_;
 wire _2622_;
 wire _2623_;
 wire _2624_;
 wire _2625_;
 wire _2626_;
 wire _2627_;
 wire _2628_;
 wire _2629_;
 wire _2630_;
 wire _2631_;
 wire _2632_;
 wire _2633_;
 wire _2634_;
 wire _2635_;
 wire _2636_;
 wire _2637_;
 wire _2638_;
 wire _2639_;
 wire _2640_;
 wire _2641_;
 wire _2642_;
 wire _2643_;
 wire _2644_;
 wire _2645_;
 wire _2646_;
 wire _2647_;
 wire _2648_;
 wire _2649_;
 wire _2650_;
 wire _2651_;
 wire _2652_;
 wire _2653_;
 wire _2654_;
 wire _2655_;
 wire _2656_;
 wire _2657_;
 wire _2658_;
 wire _2659_;
 wire _2660_;
 wire _2661_;
 wire _2662_;
 wire _2663_;
 wire _2664_;
 wire _2665_;
 wire _2666_;
 wire _2667_;
 wire _2668_;
 wire _2669_;
 wire _2670_;
 wire _2671_;
 wire _2672_;
 wire _2673_;
 wire _2674_;
 wire _2675_;
 wire _2676_;
 wire _2677_;
 wire _2678_;
 wire _2679_;
 wire _2680_;
 wire _2681_;
 wire _2682_;
 wire _2683_;
 wire _2684_;
 wire _2685_;
 wire _2686_;
 wire _2687_;
 wire _2688_;
 wire _2689_;
 wire _2690_;
 wire _2691_;
 wire _2692_;
 wire _2693_;
 wire _2694_;
 wire _2695_;
 wire _2696_;
 wire _2697_;
 wire _2698_;
 wire _2699_;
 wire _2700_;
 wire _2701_;
 wire _2702_;
 wire _2703_;
 wire _2704_;
 wire _2705_;
 wire _2706_;
 wire _2707_;
 wire _2708_;
 wire _2709_;
 wire _2710_;
 wire _2711_;
 wire _2712_;
 wire _2713_;
 wire _2714_;
 wire _2715_;
 wire _2716_;
 wire _2717_;
 wire _2718_;
 wire _2719_;
 wire _2720_;
 wire _2721_;
 wire _2722_;
 wire _2723_;
 wire _2724_;
 wire _2725_;
 wire _2726_;
 wire _2727_;
 wire _2728_;
 wire _2729_;
 wire _2730_;
 wire _2731_;
 wire _2732_;
 wire _2733_;
 wire _2734_;
 wire _2735_;
 wire _2736_;
 wire _2737_;
 wire _2738_;
 wire _2739_;
 wire _2740_;
 wire _2741_;
 wire _2742_;
 wire _2743_;
 wire _2744_;
 wire _2745_;
 wire _2746_;
 wire _2747_;
 wire _2748_;
 wire _2749_;
 wire _2750_;
 wire _2751_;
 wire _2752_;
 wire _2753_;
 wire _2754_;
 wire _2755_;
 wire _2756_;
 wire _2757_;
 wire _2758_;
 wire _2759_;
 wire _2760_;
 wire _2761_;
 wire _2762_;
 wire _2763_;
 wire _2764_;
 wire _2765_;
 wire _2766_;
 wire _2767_;
 wire _2768_;
 wire _2769_;
 wire _2770_;
 wire _2771_;
 wire _2772_;
 wire _2773_;
 wire _2774_;
 wire _2775_;
 wire _2776_;
 wire _2777_;
 wire _2778_;
 wire _2779_;
 wire _2780_;
 wire _2781_;
 wire _2782_;
 wire _2783_;
 wire _2784_;
 wire _2785_;
 wire _2786_;
 wire _2787_;
 wire _2788_;
 wire _2789_;
 wire _2790_;
 wire _2791_;
 wire _2792_;
 wire _2793_;
 wire _2794_;
 wire _2795_;
 wire _2796_;
 wire _2797_;
 wire _2798_;
 wire _2799_;
 wire _2800_;
 wire _2801_;
 wire _2802_;
 wire _2803_;
 wire _2804_;
 wire _2805_;
 wire _2806_;
 wire _2807_;
 wire _2808_;
 wire _2809_;
 wire _2810_;
 wire _2811_;
 wire _2812_;
 wire _2813_;
 wire _2814_;
 wire _2815_;
 wire _2816_;
 wire _2817_;
 wire _2818_;
 wire _2819_;
 wire _2820_;
 wire _2821_;
 wire _2822_;
 wire _2823_;
 wire _2824_;
 wire _2825_;
 wire _2826_;
 wire _2827_;
 wire _2828_;
 wire _2829_;
 wire _2830_;
 wire _2831_;
 wire _2832_;
 wire _2833_;
 wire _2834_;
 wire _2835_;
 wire _2836_;
 wire _2837_;
 wire _2838_;
 wire _2839_;
 wire _2840_;
 wire _2841_;
 wire _2842_;
 wire _2843_;
 wire _2844_;
 wire _2845_;
 wire _2846_;
 wire _2847_;
 wire _2848_;
 wire _2849_;
 wire _2850_;
 wire _2851_;
 wire _2852_;
 wire _2853_;
 wire _2854_;
 wire _2855_;
 wire _2856_;
 wire _2857_;
 wire _2858_;
 wire _2859_;
 wire _2860_;
 wire _2861_;
 wire _2862_;
 wire _2863_;
 wire _2864_;
 wire _2865_;
 wire _2866_;
 wire _2867_;
 wire _2868_;
 wire _2869_;
 wire _2870_;
 wire _2871_;
 wire _2872_;
 wire _2873_;
 wire _2874_;
 wire _2875_;
 wire _2876_;
 wire _2877_;
 wire _2878_;
 wire _2879_;
 wire _2880_;
 wire _2881_;
 wire _2882_;
 wire _2883_;
 wire _2884_;
 wire _2885_;
 wire _2886_;
 wire _2887_;
 wire _2888_;
 wire _2889_;
 wire _2890_;
 wire _2891_;
 wire _2892_;
 wire _2893_;
 wire _2894_;
 wire _2895_;
 wire _2896_;
 wire _2897_;
 wire _2898_;
 wire _2899_;
 wire _2900_;
 wire _2901_;
 wire _2902_;
 wire _2903_;
 wire _2904_;
 wire _2905_;
 wire _2906_;
 wire _2907_;
 wire _2908_;
 wire _2909_;
 wire _2910_;
 wire _2911_;
 wire _2912_;
 wire _2913_;
 wire _2914_;
 wire _2915_;
 wire _2916_;
 wire _2917_;
 wire _2918_;
 wire _2919_;
 wire _2920_;
 wire _2921_;
 wire _2922_;
 wire _2923_;
 wire _2924_;
 wire _2925_;
 wire _2926_;
 wire _2927_;
 wire _2928_;
 wire _2929_;
 wire _2930_;
 wire _2931_;
 wire _2932_;
 wire _2933_;
 wire _2934_;
 wire _2935_;
 wire _2936_;
 wire _2937_;
 wire _2938_;
 wire _2939_;
 wire _2940_;
 wire _2941_;
 wire _2942_;
 wire _2943_;
 wire _2944_;
 wire _2945_;
 wire _2946_;
 wire _2947_;
 wire _2948_;
 wire _2949_;
 wire _2950_;
 wire _2951_;
 wire _2952_;
 wire _2953_;
 wire _2954_;
 wire _2955_;
 wire _2956_;
 wire _2957_;
 wire _2958_;
 wire _2959_;
 wire _2960_;
 wire _2961_;
 wire _2962_;
 wire _2963_;
 wire _2964_;
 wire _2965_;
 wire _2966_;
 wire _2967_;
 wire _2968_;
 wire _2969_;
 wire _2970_;
 wire _2971_;
 wire _2972_;
 wire _2973_;
 wire _2974_;
 wire _2975_;
 wire _2976_;
 wire _2977_;
 wire _2978_;
 wire _2979_;
 wire _2980_;
 wire _2981_;
 wire _2982_;
 wire _2983_;
 wire _2984_;
 wire _2985_;
 wire _2986_;
 wire _2987_;
 wire _2988_;
 wire _2989_;
 wire _2990_;
 wire _2991_;
 wire _2992_;
 wire _2993_;
 wire _2994_;
 wire _2995_;
 wire _2996_;
 wire _2997_;
 wire _2998_;
 wire _2999_;
 wire _3000_;
 wire _3001_;
 wire _3002_;
 wire _3003_;
 wire _3004_;
 wire _3005_;
 wire _3006_;
 wire _3007_;
 wire _3008_;
 wire _3009_;
 wire _3010_;
 wire _3011_;
 wire _3012_;
 wire _3013_;
 wire _3014_;
 wire _3015_;
 wire _3016_;
 wire _3017_;
 wire _3018_;
 wire _3019_;
 wire _3020_;
 wire _3021_;
 wire _3022_;
 wire _3023_;
 wire _3024_;
 wire _3025_;
 wire _3026_;
 wire _3027_;
 wire _3028_;
 wire _3029_;
 wire _3030_;
 wire _3031_;
 wire _3032_;
 wire _3033_;
 wire _3034_;
 wire _3035_;
 wire _3036_;
 wire _3037_;
 wire _3038_;
 wire _3039_;
 wire _3040_;
 wire _3041_;
 wire _3042_;
 wire _3043_;
 wire _3044_;
 wire _3045_;
 wire _3046_;
 wire _3047_;
 wire _3048_;
 wire _3049_;
 wire _3050_;
 wire _3051_;
 wire _3052_;
 wire _3053_;
 wire _3054_;
 wire _3055_;
 wire _3056_;
 wire _3057_;
 wire _3058_;
 wire _3059_;
 wire _3060_;
 wire _3061_;
 wire _3062_;
 wire _3063_;
 wire _3064_;
 wire _3065_;
 wire _3066_;
 wire _3067_;
 wire _3068_;
 wire _3069_;
 wire _3070_;
 wire _3071_;
 wire _3072_;
 wire _3073_;
 wire _3074_;
 wire _3075_;
 wire _3076_;
 wire _3077_;
 wire _3078_;
 wire _3079_;
 wire _3080_;
 wire _3081_;
 wire _3082_;
 wire _3083_;
 wire _3084_;
 wire _3085_;
 wire _3086_;
 wire _3087_;
 wire _3088_;
 wire _3089_;
 wire _3090_;
 wire _3091_;
 wire _3092_;
 wire _3093_;
 wire _3094_;
 wire _3095_;
 wire _3096_;
 wire _3097_;
 wire _3098_;
 wire _3099_;
 wire _3100_;
 wire _3101_;
 wire _3102_;
 wire _3103_;
 wire _3104_;
 wire _3105_;
 wire _3106_;
 wire _3107_;
 wire _3108_;
 wire _3109_;
 wire _3110_;
 wire _3111_;
 wire _3112_;
 wire _3113_;
 wire _3114_;
 wire _3115_;
 wire _3116_;
 wire _3117_;
 wire _3118_;
 wire _3119_;
 wire _3120_;
 wire _3121_;
 wire _3122_;
 wire _3123_;
 wire _3124_;
 wire _3125_;
 wire _3126_;
 wire _3127_;
 wire _3128_;
 wire _3129_;
 wire _3130_;
 wire _3131_;
 wire _3132_;
 wire _3133_;
 wire _3134_;
 wire _3135_;
 wire _3136_;
 wire _3137_;
 wire _3138_;
 wire _3139_;
 wire _3140_;
 wire _3141_;
 wire _3142_;
 wire _3143_;
 wire _3144_;
 wire _3145_;
 wire _3146_;
 wire _3147_;
 wire _3148_;
 wire _3149_;
 wire _3150_;
 wire _3151_;
 wire _3152_;
 wire _3153_;
 wire _3154_;
 wire _3155_;
 wire _3156_;
 wire _3157_;
 wire _3158_;
 wire _3159_;
 wire _3160_;
 wire _3161_;
 wire _3162_;
 wire _3163_;
 wire _3164_;
 wire _3165_;
 wire _3166_;
 wire _3167_;
 wire _3168_;
 wire _3169_;
 wire _3170_;
 wire _3171_;
 wire _3172_;
 wire _3173_;
 wire _3174_;
 wire _3175_;
 wire _3176_;
 wire _3177_;
 wire _3178_;
 wire _3179_;
 wire _3180_;
 wire _3181_;
 wire _3182_;
 wire _3183_;
 wire _3184_;
 wire _3185_;
 wire _3186_;
 wire _3187_;
 wire _3188_;
 wire _3189_;
 wire _3190_;
 wire _3191_;
 wire _3192_;
 wire _3193_;
 wire _3194_;
 wire _3195_;
 wire _3196_;
 wire _3197_;
 wire _3198_;
 wire _3199_;
 wire _3200_;
 wire _3201_;
 wire _3202_;
 wire _3203_;
 wire _3204_;
 wire _3205_;
 wire _3206_;
 wire _3207_;
 wire _3208_;
 wire _3209_;
 wire _3210_;
 wire _3211_;
 wire _3212_;
 wire _3213_;
 wire _3214_;
 wire _3215_;
 wire _3216_;
 wire _3217_;
 wire _3218_;
 wire _3219_;
 wire _3220_;
 wire _3221_;
 wire _3222_;
 wire _3223_;
 wire _3224_;
 wire _3225_;
 wire _3226_;
 wire _3227_;
 wire _3228_;
 wire _3229_;
 wire _3230_;
 wire _3231_;
 wire _3232_;
 wire _3233_;
 wire _3234_;
 wire _3235_;
 wire _3236_;
 wire _3237_;
 wire _3238_;
 wire _3239_;
 wire _3240_;
 wire _3241_;
 wire _3242_;
 wire _3243_;
 wire _3244_;
 wire _3245_;
 wire _3246_;
 wire _3247_;
 wire _3248_;
 wire _3249_;
 wire _3250_;
 wire _3251_;
 wire _3252_;
 wire _3253_;
 wire _3254_;
 wire _3255_;
 wire _3256_;
 wire _3257_;
 wire _3258_;
 wire _3259_;
 wire _3260_;
 wire _3261_;
 wire _3262_;
 wire _3263_;
 wire _3264_;
 wire _3265_;
 wire _3266_;
 wire _3267_;
 wire _3268_;
 wire _3269_;
 wire _3270_;
 wire _3271_;
 wire _3272_;
 wire _3273_;
 wire _3274_;
 wire _3275_;
 wire _3276_;
 wire _3277_;
 wire _3278_;
 wire _3279_;
 wire _3280_;
 wire _3281_;
 wire _3282_;
 wire _3283_;
 wire _3284_;
 wire _3285_;
 wire _3286_;
 wire _3287_;
 wire _3288_;
 wire _3289_;
 wire _3290_;
 wire _3291_;
 wire _3292_;
 wire _3293_;
 wire _3294_;
 wire _3295_;
 wire _3296_;
 wire _3297_;
 wire _3298_;
 wire _3299_;
 wire _3300_;
 wire _3301_;
 wire _3302_;
 wire _3303_;
 wire _3304_;
 wire _3305_;
 wire _3306_;
 wire _3307_;
 wire _3308_;
 wire _3309_;
 wire _3310_;
 wire _3311_;
 wire _3312_;
 wire _3313_;
 wire _3314_;
 wire _3315_;
 wire _3316_;
 wire _3317_;
 wire _3318_;
 wire _3319_;
 wire _3320_;
 wire _3321_;
 wire _3322_;
 wire _3323_;
 wire _3324_;
 wire _3325_;
 wire _3326_;
 wire _3327_;
 wire _3328_;
 wire _3329_;
 wire _3330_;
 wire _3331_;
 wire _3332_;
 wire _3333_;
 wire _3334_;
 wire _3335_;
 wire _3336_;
 wire _3337_;
 wire _3338_;
 wire _3339_;
 wire _3340_;
 wire _3341_;
 wire _3342_;
 wire _3343_;
 wire _3344_;
 wire _3345_;
 wire _3346_;
 wire _3347_;
 wire _3348_;
 wire _3349_;
 wire _3350_;
 wire _3351_;
 wire _3352_;
 wire _3353_;
 wire _3354_;
 wire _3355_;
 wire _3356_;
 wire _3357_;
 wire _3358_;
 wire _3359_;
 wire _3360_;
 wire _3361_;
 wire _3362_;
 wire _3363_;
 wire _3364_;
 wire _3365_;
 wire _3366_;
 wire _3367_;
 wire _3368_;
 wire _3369_;
 wire _3370_;
 wire _3371_;
 wire _3372_;
 wire _3373_;
 wire _3374_;
 wire _3375_;
 wire _3376_;
 wire _3377_;
 wire _3378_;
 wire _3379_;
 wire _3380_;
 wire _3381_;
 wire _3382_;
 wire _3383_;
 wire _3384_;
 wire _3385_;
 wire _3386_;
 wire _3387_;
 wire _3388_;
 wire _3389_;
 wire _3390_;
 wire _3391_;
 wire _3392_;
 wire _3393_;
 wire _3394_;
 wire _3395_;
 wire _3396_;
 wire _3397_;
 wire _3398_;
 wire _3399_;
 wire _3400_;
 wire _3401_;
 wire _3402_;
 wire _3403_;
 wire _3404_;
 wire _3405_;
 wire _3406_;
 wire _3407_;
 wire _3408_;
 wire _3409_;
 wire _3410_;
 wire _3411_;
 wire _3412_;
 wire _3413_;
 wire _3414_;
 wire _3415_;
 wire _3416_;
 wire _3417_;
 wire _3418_;
 wire _3419_;
 wire _3420_;
 wire _3421_;
 wire _3422_;
 wire _3423_;
 wire _3424_;
 wire _3425_;
 wire _3426_;
 wire _3427_;
 wire _3428_;
 wire _3429_;
 wire _3430_;
 wire _3431_;
 wire _3432_;
 wire _3433_;
 wire _3434_;
 wire _3435_;
 wire _3436_;
 wire _3437_;
 wire _3438_;
 wire _3439_;
 wire _3440_;
 wire _3441_;
 wire _3442_;
 wire _3443_;
 wire _3444_;
 wire _3445_;
 wire _3446_;
 wire _3447_;
 wire _3448_;
 wire _3449_;
 wire _3450_;
 wire _3451_;
 wire _3452_;
 wire _3453_;
 wire _3454_;
 wire _3455_;
 wire _3456_;
 wire _3457_;
 wire _3458_;
 wire _3459_;
 wire _3460_;
 wire _3461_;
 wire _3462_;
 wire _3463_;
 wire _3464_;
 wire _3465_;
 wire _3466_;
 wire _3467_;
 wire _3468_;
 wire _3469_;
 wire _3470_;
 wire _3471_;
 wire _3472_;
 wire _3473_;
 wire _3474_;
 wire _3475_;
 wire _3476_;
 wire _3477_;
 wire _3478_;
 wire _3479_;
 wire _3480_;
 wire _3481_;
 wire _3482_;
 wire _3483_;
 wire _3484_;
 wire _3485_;
 wire _3486_;
 wire _3487_;
 wire _3488_;
 wire _3489_;
 wire _3490_;
 wire _3491_;
 wire _3492_;
 wire _3493_;
 wire _3494_;
 wire _3495_;
 wire _3496_;
 wire _3497_;
 wire _3498_;
 wire _3499_;
 wire _3500_;
 wire _3501_;
 wire _3502_;
 wire _3503_;
 wire _3504_;
 wire _3505_;
 wire _3506_;
 wire _3507_;
 wire _3508_;
 wire _3509_;
 wire _3510_;
 wire _3511_;
 wire _3512_;
 wire _3513_;
 wire _3514_;
 wire _3515_;
 wire _3516_;
 wire _3517_;
 wire _3518_;
 wire _3519_;
 wire _3520_;
 wire _3521_;
 wire _3522_;
 wire _3523_;
 wire _3524_;
 wire _3525_;
 wire _3526_;
 wire _3527_;
 wire _3528_;
 wire _3529_;
 wire _3530_;
 wire _3531_;
 wire _3532_;
 wire _3533_;
 wire _3534_;
 wire _3535_;
 wire _3536_;
 wire _3537_;
 wire _3538_;
 wire _3539_;
 wire _3540_;
 wire _3541_;
 wire _3542_;
 wire _3543_;
 wire _3544_;
 wire _3545_;
 wire _3546_;
 wire _3547_;
 wire _3548_;
 wire _3549_;
 wire _3550_;
 wire _3551_;
 wire _3552_;
 wire _3553_;
 wire _3554_;
 wire _3555_;
 wire _3556_;
 wire _3557_;
 wire _3558_;
 wire _3559_;
 wire _3560_;
 wire _3561_;
 wire _3562_;
 wire _3563_;
 wire _3564_;
 wire _3565_;
 wire _3566_;
 wire _3567_;
 wire _3568_;
 wire _3569_;
 wire _3570_;
 wire _3571_;
 wire _3572_;
 wire _3573_;
 wire _3574_;
 wire _3575_;
 wire _3576_;
 wire _3577_;
 wire _3578_;
 wire _3579_;
 wire _3580_;
 wire _3581_;
 wire _3582_;
 wire _3583_;
 wire _3584_;
 wire _3585_;
 wire _3586_;
 wire _3587_;
 wire _3588_;
 wire _3589_;
 wire _3590_;
 wire _3591_;
 wire _3592_;
 wire _3593_;
 wire _3594_;
 wire _3595_;
 wire _3596_;
 wire _3597_;
 wire _3598_;
 wire _3599_;
 wire _3600_;
 wire _3601_;
 wire _3602_;
 wire _3603_;
 wire _3604_;
 wire _3605_;
 wire _3606_;
 wire _3607_;
 wire _3608_;
 wire _3609_;
 wire _3610_;
 wire _3611_;
 wire _3612_;
 wire _3613_;
 wire _3614_;
 wire _3615_;
 wire _3616_;
 wire _3617_;
 wire _3618_;
 wire _3619_;
 wire _3620_;
 wire _3621_;
 wire _3622_;
 wire _3623_;
 wire _3624_;
 wire _3625_;
 wire _3626_;
 wire _3627_;
 wire _3628_;
 wire _3629_;
 wire _3630_;
 wire _3631_;
 wire _3632_;
 wire _3633_;
 wire _3634_;
 wire _3635_;
 wire _3636_;
 wire _3637_;
 wire _3638_;
 wire _3639_;
 wire _3640_;
 wire _3641_;
 wire _3642_;
 wire _3643_;
 wire _3644_;
 wire _3645_;
 wire _3646_;
 wire _3647_;
 wire _3648_;
 wire _3649_;
 wire _3650_;
 wire _3651_;
 wire _3652_;
 wire _3653_;
 wire _3654_;
 wire _3655_;
 wire _3656_;
 wire _3657_;
 wire _3658_;
 wire _3659_;
 wire _3660_;
 wire _3661_;
 wire _3662_;
 wire _3663_;
 wire _3664_;
 wire _3665_;
 wire _3666_;
 wire _3667_;
 wire _3668_;
 wire _3669_;
 wire _3670_;
 wire _3671_;
 wire _3672_;
 wire _3673_;
 wire _3674_;
 wire _3675_;
 wire _3676_;
 wire _3677_;
 wire _3678_;
 wire _3679_;
 wire _3680_;
 wire _3681_;
 wire _3682_;
 wire _3683_;
 wire _3684_;
 wire _3685_;
 wire _3686_;
 wire _3687_;
 wire _3688_;
 wire _3689_;
 wire _3690_;
 wire _3691_;
 wire _3692_;
 wire _3693_;
 wire _3694_;
 wire _3695_;
 wire _3696_;
 wire _3697_;
 wire _3698_;
 wire _3699_;
 wire _3700_;
 wire _3701_;
 wire _3702_;
 wire _3703_;
 wire _3704_;
 wire _3705_;
 wire _3706_;
 wire _3707_;
 wire _3708_;
 wire _3709_;
 wire _3710_;
 wire _3711_;
 wire _3712_;
 wire _3713_;
 wire _3714_;
 wire _3715_;
 wire _3716_;
 wire _3717_;
 wire _3718_;
 wire _3719_;
 wire _3720_;
 wire _3721_;
 wire _3722_;
 wire _3723_;
 wire _3724_;
 wire _3725_;
 wire _3726_;
 wire _3727_;
 wire _3728_;
 wire _3729_;
 wire _3730_;
 wire _3731_;
 wire _3732_;
 wire _3733_;
 wire _3734_;
 wire _3735_;
 wire _3736_;
 wire _3737_;
 wire _3738_;
 wire _3739_;
 wire _3740_;
 wire _3741_;
 wire _3742_;
 wire _3743_;
 wire _3744_;
 wire _3745_;
 wire _3746_;
 wire _3747_;
 wire _3748_;
 wire _3749_;
 wire _3750_;
 wire _3751_;
 wire _3752_;
 wire _3753_;
 wire _3754_;
 wire _3755_;
 wire _3756_;
 wire _3757_;
 wire _3758_;
 wire _3759_;
 wire _3760_;
 wire _3761_;
 wire _3762_;
 wire _3763_;
 wire _3764_;
 wire _3765_;
 wire _3766_;
 wire _3767_;
 wire _3768_;
 wire _3769_;
 wire _3770_;
 wire _3771_;
 wire _3772_;
 wire _3773_;
 wire _3774_;
 wire _3775_;
 wire _3776_;
 wire _3777_;
 wire _3778_;
 wire _3779_;
 wire _3780_;
 wire _3781_;
 wire _3782_;
 wire _3783_;
 wire _3784_;
 wire _3785_;
 wire _3786_;
 wire _3787_;
 wire _3788_;
 wire _3789_;
 wire _3790_;
 wire _3791_;
 wire _3792_;
 wire _3793_;
 wire _3794_;
 wire _3795_;
 wire _3796_;
 wire _3797_;
 wire _3798_;
 wire _3799_;
 wire _3800_;
 wire _3801_;
 wire _3802_;
 wire _3803_;
 wire _3804_;
 wire _3805_;
 wire _3806_;
 wire _3807_;
 wire _3808_;
 wire _3809_;
 wire _3810_;
 wire _3811_;
 wire _3812_;
 wire _3813_;
 wire _3814_;
 wire _3815_;
 wire _3816_;
 wire _3817_;
 wire _3818_;
 wire _3819_;
 wire _3820_;
 wire _3821_;
 wire _3822_;
 wire _3823_;
 wire _3824_;
 wire _3825_;
 wire _3826_;
 wire _3827_;
 wire _3828_;
 wire _3829_;
 wire _3830_;
 wire _3831_;
 wire _3832_;
 wire _3833_;
 wire _3834_;
 wire _3835_;
 wire _3836_;
 wire _3837_;
 wire _3838_;
 wire _3839_;
 wire _3840_;
 wire _3841_;
 wire _3842_;
 wire _3843_;
 wire _3844_;
 wire _3845_;
 wire _3846_;
 wire _3847_;
 wire _3848_;
 wire _3849_;
 wire _3850_;
 wire _3851_;
 wire _3852_;
 wire _3853_;
 wire _3854_;
 wire _3855_;
 wire _3856_;
 wire _3857_;
 wire _3858_;
 wire _3859_;
 wire _3860_;
 wire _3861_;
 wire _3862_;
 wire _3863_;
 wire _3864_;
 wire _3865_;
 wire _3866_;
 wire _3867_;
 wire _3868_;
 wire _3869_;
 wire _3870_;
 wire _3871_;
 wire _3872_;
 wire _3873_;
 wire _3874_;
 wire _3875_;
 wire _3876_;
 wire _3877_;
 wire _3878_;
 wire _3879_;
 wire _3880_;
 wire _3881_;
 wire _3882_;
 wire _3883_;
 wire _3884_;
 wire _3885_;
 wire _3886_;
 wire _3887_;
 wire _3888_;
 wire _3889_;
 wire _3890_;
 wire _3891_;
 wire _3892_;
 wire _3893_;
 wire _3894_;
 wire _3895_;
 wire _3896_;
 wire _3897_;
 wire _3898_;
 wire _3899_;
 wire _3900_;
 wire _3901_;
 wire _3902_;
 wire _3903_;
 wire _3904_;
 wire _3905_;
 wire _3906_;
 wire _3907_;
 wire _3908_;
 wire _3909_;
 wire _3910_;
 wire _3911_;
 wire _3912_;
 wire _3913_;
 wire _3914_;
 wire _3915_;
 wire _3916_;
 wire _3917_;
 wire _3918_;
 wire _3919_;
 wire _3920_;
 wire _3921_;
 wire _3922_;
 wire _3923_;
 wire _3924_;
 wire _3925_;
 wire _3926_;
 wire _3927_;
 wire _3928_;
 wire _3929_;
 wire _3930_;
 wire _3931_;
 wire net12;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net13;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net14;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net50;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net51;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net52;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net80;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net81;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net82;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net83;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net84;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net85;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire \mod.Arithmetic.ACTI.x[0] ;
 wire \mod.Arithmetic.ACTI.x[1] ;
 wire \mod.Arithmetic.ACTI.x[2] ;
 wire \mod.Arithmetic.ACTI.x[3] ;
 wire \mod.Arithmetic.ACTI.x[4] ;
 wire \mod.Arithmetic.ACTI.x[5] ;
 wire \mod.Arithmetic.ACTI.x[6] ;
 wire \mod.Arithmetic.ACTI.x[7] ;
 wire \mod.Arithmetic.CN.F_in[0] ;
 wire \mod.Arithmetic.CN.I_in[10] ;
 wire \mod.Arithmetic.CN.I_in[11] ;
 wire \mod.Arithmetic.CN.I_in[12] ;
 wire \mod.Arithmetic.CN.I_in[13] ;
 wire \mod.Arithmetic.CN.I_in[14] ;
 wire \mod.Arithmetic.CN.I_in[15] ;
 wire \mod.Arithmetic.CN.I_in[16] ;
 wire \mod.Arithmetic.CN.I_in[17] ;
 wire \mod.Arithmetic.CN.I_in[18] ;
 wire \mod.Arithmetic.CN.I_in[19] ;
 wire \mod.Arithmetic.CN.I_in[20] ;
 wire \mod.Arithmetic.CN.I_in[21] ;
 wire \mod.Arithmetic.CN.I_in[22] ;
 wire \mod.Arithmetic.CN.I_in[23] ;
 wire \mod.Arithmetic.CN.I_in[24] ;
 wire \mod.Arithmetic.CN.I_in[25] ;
 wire \mod.Arithmetic.CN.I_in[26] ;
 wire \mod.Arithmetic.CN.I_in[27] ;
 wire \mod.Arithmetic.CN.I_in[28] ;
 wire \mod.Arithmetic.CN.I_in[29] ;
 wire \mod.Arithmetic.CN.I_in[30] ;
 wire \mod.Arithmetic.CN.I_in[31] ;
 wire \mod.Arithmetic.CN.I_in[32] ;
 wire \mod.Arithmetic.CN.I_in[33] ;
 wire \mod.Arithmetic.CN.I_in[34] ;
 wire \mod.Arithmetic.CN.I_in[35] ;
 wire \mod.Arithmetic.CN.I_in[36] ;
 wire \mod.Arithmetic.CN.I_in[37] ;
 wire \mod.Arithmetic.CN.I_in[38] ;
 wire \mod.Arithmetic.CN.I_in[39] ;
 wire \mod.Arithmetic.CN.I_in[40] ;
 wire \mod.Arithmetic.CN.I_in[41] ;
 wire \mod.Arithmetic.CN.I_in[42] ;
 wire \mod.Arithmetic.CN.I_in[43] ;
 wire \mod.Arithmetic.CN.I_in[44] ;
 wire \mod.Arithmetic.CN.I_in[45] ;
 wire \mod.Arithmetic.CN.I_in[46] ;
 wire \mod.Arithmetic.CN.I_in[47] ;
 wire \mod.Arithmetic.CN.I_in[48] ;
 wire \mod.Arithmetic.CN.I_in[49] ;
 wire \mod.Arithmetic.CN.I_in[50] ;
 wire \mod.Arithmetic.CN.I_in[51] ;
 wire \mod.Arithmetic.CN.I_in[52] ;
 wire \mod.Arithmetic.CN.I_in[53] ;
 wire \mod.Arithmetic.CN.I_in[54] ;
 wire \mod.Arithmetic.CN.I_in[55] ;
 wire \mod.Arithmetic.CN.I_in[56] ;
 wire \mod.Arithmetic.CN.I_in[57] ;
 wire \mod.Arithmetic.CN.I_in[58] ;
 wire \mod.Arithmetic.CN.I_in[59] ;
 wire \mod.Arithmetic.CN.I_in[60] ;
 wire \mod.Arithmetic.CN.I_in[61] ;
 wire \mod.Arithmetic.CN.I_in[62] ;
 wire \mod.Arithmetic.CN.I_in[63] ;
 wire \mod.Arithmetic.CN.I_in[64] ;
 wire \mod.Arithmetic.CN.I_in[65] ;
 wire \mod.Arithmetic.CN.I_in[66] ;
 wire \mod.Arithmetic.CN.I_in[67] ;
 wire \mod.Arithmetic.CN.I_in[68] ;
 wire \mod.Arithmetic.CN.I_in[69] ;
 wire \mod.Arithmetic.CN.I_in[70] ;
 wire \mod.Arithmetic.CN.I_in[71] ;
 wire \mod.Arithmetic.CN.I_in[8] ;
 wire \mod.Arithmetic.CN.I_in[9] ;
 wire \mod.Arithmetic.I_out[72] ;
 wire \mod.Arithmetic.I_out[73] ;
 wire \mod.Arithmetic.I_out[74] ;
 wire \mod.Arithmetic.I_out[75] ;
 wire \mod.Arithmetic.I_out[76] ;
 wire \mod.Arithmetic.I_out[77] ;
 wire \mod.Arithmetic.I_out[78] ;
 wire \mod.Arithmetic.I_out[79] ;
 wire \mod.DM_en ;
 wire \mod.DMen_reg ;
 wire \mod.DMen_reg2 ;
 wire \mod.Data_Mem.F_M.MRAM[0][0] ;
 wire \mod.Data_Mem.F_M.MRAM[0][1] ;
 wire \mod.Data_Mem.F_M.MRAM[0][2] ;
 wire \mod.Data_Mem.F_M.MRAM[0][3] ;
 wire \mod.Data_Mem.F_M.MRAM[0][4] ;
 wire \mod.Data_Mem.F_M.MRAM[0][5] ;
 wire \mod.Data_Mem.F_M.MRAM[0][6] ;
 wire \mod.Data_Mem.F_M.MRAM[0][7] ;
 wire \mod.Data_Mem.F_M.MRAM[10][0] ;
 wire \mod.Data_Mem.F_M.MRAM[10][1] ;
 wire \mod.Data_Mem.F_M.MRAM[10][2] ;
 wire \mod.Data_Mem.F_M.MRAM[10][3] ;
 wire \mod.Data_Mem.F_M.MRAM[10][4] ;
 wire \mod.Data_Mem.F_M.MRAM[10][5] ;
 wire \mod.Data_Mem.F_M.MRAM[10][6] ;
 wire \mod.Data_Mem.F_M.MRAM[10][7] ;
 wire \mod.Data_Mem.F_M.MRAM[11][0] ;
 wire \mod.Data_Mem.F_M.MRAM[11][1] ;
 wire \mod.Data_Mem.F_M.MRAM[11][2] ;
 wire \mod.Data_Mem.F_M.MRAM[11][3] ;
 wire \mod.Data_Mem.F_M.MRAM[11][4] ;
 wire \mod.Data_Mem.F_M.MRAM[11][5] ;
 wire \mod.Data_Mem.F_M.MRAM[11][6] ;
 wire \mod.Data_Mem.F_M.MRAM[11][7] ;
 wire \mod.Data_Mem.F_M.MRAM[12][0] ;
 wire \mod.Data_Mem.F_M.MRAM[12][1] ;
 wire \mod.Data_Mem.F_M.MRAM[12][2] ;
 wire \mod.Data_Mem.F_M.MRAM[12][3] ;
 wire \mod.Data_Mem.F_M.MRAM[12][4] ;
 wire \mod.Data_Mem.F_M.MRAM[12][5] ;
 wire \mod.Data_Mem.F_M.MRAM[12][6] ;
 wire \mod.Data_Mem.F_M.MRAM[12][7] ;
 wire \mod.Data_Mem.F_M.MRAM[13][0] ;
 wire \mod.Data_Mem.F_M.MRAM[13][1] ;
 wire \mod.Data_Mem.F_M.MRAM[13][2] ;
 wire \mod.Data_Mem.F_M.MRAM[13][3] ;
 wire \mod.Data_Mem.F_M.MRAM[13][4] ;
 wire \mod.Data_Mem.F_M.MRAM[13][5] ;
 wire \mod.Data_Mem.F_M.MRAM[13][6] ;
 wire \mod.Data_Mem.F_M.MRAM[13][7] ;
 wire \mod.Data_Mem.F_M.MRAM[14][0] ;
 wire \mod.Data_Mem.F_M.MRAM[14][1] ;
 wire \mod.Data_Mem.F_M.MRAM[14][2] ;
 wire \mod.Data_Mem.F_M.MRAM[14][3] ;
 wire \mod.Data_Mem.F_M.MRAM[14][4] ;
 wire \mod.Data_Mem.F_M.MRAM[14][5] ;
 wire \mod.Data_Mem.F_M.MRAM[14][6] ;
 wire \mod.Data_Mem.F_M.MRAM[14][7] ;
 wire \mod.Data_Mem.F_M.MRAM[15][0] ;
 wire \mod.Data_Mem.F_M.MRAM[15][1] ;
 wire \mod.Data_Mem.F_M.MRAM[15][2] ;
 wire \mod.Data_Mem.F_M.MRAM[15][3] ;
 wire \mod.Data_Mem.F_M.MRAM[15][4] ;
 wire \mod.Data_Mem.F_M.MRAM[15][5] ;
 wire \mod.Data_Mem.F_M.MRAM[15][6] ;
 wire \mod.Data_Mem.F_M.MRAM[15][7] ;
 wire \mod.Data_Mem.F_M.MRAM[16][0] ;
 wire \mod.Data_Mem.F_M.MRAM[16][1] ;
 wire \mod.Data_Mem.F_M.MRAM[16][2] ;
 wire \mod.Data_Mem.F_M.MRAM[16][3] ;
 wire \mod.Data_Mem.F_M.MRAM[16][4] ;
 wire \mod.Data_Mem.F_M.MRAM[16][5] ;
 wire \mod.Data_Mem.F_M.MRAM[16][6] ;
 wire \mod.Data_Mem.F_M.MRAM[16][7] ;
 wire \mod.Data_Mem.F_M.MRAM[17][0] ;
 wire \mod.Data_Mem.F_M.MRAM[17][1] ;
 wire \mod.Data_Mem.F_M.MRAM[17][2] ;
 wire \mod.Data_Mem.F_M.MRAM[17][3] ;
 wire \mod.Data_Mem.F_M.MRAM[17][4] ;
 wire \mod.Data_Mem.F_M.MRAM[17][5] ;
 wire \mod.Data_Mem.F_M.MRAM[17][6] ;
 wire \mod.Data_Mem.F_M.MRAM[17][7] ;
 wire \mod.Data_Mem.F_M.MRAM[18][0] ;
 wire \mod.Data_Mem.F_M.MRAM[18][1] ;
 wire \mod.Data_Mem.F_M.MRAM[18][2] ;
 wire \mod.Data_Mem.F_M.MRAM[18][3] ;
 wire \mod.Data_Mem.F_M.MRAM[18][4] ;
 wire \mod.Data_Mem.F_M.MRAM[18][5] ;
 wire \mod.Data_Mem.F_M.MRAM[18][6] ;
 wire \mod.Data_Mem.F_M.MRAM[18][7] ;
 wire \mod.Data_Mem.F_M.MRAM[19][0] ;
 wire \mod.Data_Mem.F_M.MRAM[19][1] ;
 wire \mod.Data_Mem.F_M.MRAM[19][2] ;
 wire \mod.Data_Mem.F_M.MRAM[19][3] ;
 wire \mod.Data_Mem.F_M.MRAM[19][4] ;
 wire \mod.Data_Mem.F_M.MRAM[19][5] ;
 wire \mod.Data_Mem.F_M.MRAM[19][6] ;
 wire \mod.Data_Mem.F_M.MRAM[19][7] ;
 wire \mod.Data_Mem.F_M.MRAM[1][0] ;
 wire \mod.Data_Mem.F_M.MRAM[1][1] ;
 wire \mod.Data_Mem.F_M.MRAM[1][2] ;
 wire \mod.Data_Mem.F_M.MRAM[1][3] ;
 wire \mod.Data_Mem.F_M.MRAM[1][4] ;
 wire \mod.Data_Mem.F_M.MRAM[1][5] ;
 wire \mod.Data_Mem.F_M.MRAM[1][6] ;
 wire \mod.Data_Mem.F_M.MRAM[1][7] ;
 wire \mod.Data_Mem.F_M.MRAM[20][0] ;
 wire \mod.Data_Mem.F_M.MRAM[20][1] ;
 wire \mod.Data_Mem.F_M.MRAM[20][2] ;
 wire \mod.Data_Mem.F_M.MRAM[20][3] ;
 wire \mod.Data_Mem.F_M.MRAM[20][4] ;
 wire \mod.Data_Mem.F_M.MRAM[20][5] ;
 wire \mod.Data_Mem.F_M.MRAM[20][6] ;
 wire \mod.Data_Mem.F_M.MRAM[20][7] ;
 wire \mod.Data_Mem.F_M.MRAM[21][0] ;
 wire \mod.Data_Mem.F_M.MRAM[21][1] ;
 wire \mod.Data_Mem.F_M.MRAM[21][2] ;
 wire \mod.Data_Mem.F_M.MRAM[21][3] ;
 wire \mod.Data_Mem.F_M.MRAM[21][4] ;
 wire \mod.Data_Mem.F_M.MRAM[21][5] ;
 wire \mod.Data_Mem.F_M.MRAM[21][6] ;
 wire \mod.Data_Mem.F_M.MRAM[21][7] ;
 wire \mod.Data_Mem.F_M.MRAM[22][0] ;
 wire \mod.Data_Mem.F_M.MRAM[22][1] ;
 wire \mod.Data_Mem.F_M.MRAM[22][2] ;
 wire \mod.Data_Mem.F_M.MRAM[22][3] ;
 wire \mod.Data_Mem.F_M.MRAM[22][4] ;
 wire \mod.Data_Mem.F_M.MRAM[22][5] ;
 wire \mod.Data_Mem.F_M.MRAM[22][6] ;
 wire \mod.Data_Mem.F_M.MRAM[22][7] ;
 wire \mod.Data_Mem.F_M.MRAM[23][0] ;
 wire \mod.Data_Mem.F_M.MRAM[23][1] ;
 wire \mod.Data_Mem.F_M.MRAM[23][2] ;
 wire \mod.Data_Mem.F_M.MRAM[23][3] ;
 wire \mod.Data_Mem.F_M.MRAM[23][4] ;
 wire \mod.Data_Mem.F_M.MRAM[23][5] ;
 wire \mod.Data_Mem.F_M.MRAM[23][6] ;
 wire \mod.Data_Mem.F_M.MRAM[23][7] ;
 wire \mod.Data_Mem.F_M.MRAM[24][0] ;
 wire \mod.Data_Mem.F_M.MRAM[24][1] ;
 wire \mod.Data_Mem.F_M.MRAM[24][2] ;
 wire \mod.Data_Mem.F_M.MRAM[24][3] ;
 wire \mod.Data_Mem.F_M.MRAM[24][4] ;
 wire \mod.Data_Mem.F_M.MRAM[24][5] ;
 wire \mod.Data_Mem.F_M.MRAM[24][6] ;
 wire \mod.Data_Mem.F_M.MRAM[24][7] ;
 wire \mod.Data_Mem.F_M.MRAM[25][0] ;
 wire \mod.Data_Mem.F_M.MRAM[25][1] ;
 wire \mod.Data_Mem.F_M.MRAM[25][2] ;
 wire \mod.Data_Mem.F_M.MRAM[25][3] ;
 wire \mod.Data_Mem.F_M.MRAM[25][4] ;
 wire \mod.Data_Mem.F_M.MRAM[25][5] ;
 wire \mod.Data_Mem.F_M.MRAM[25][6] ;
 wire \mod.Data_Mem.F_M.MRAM[25][7] ;
 wire \mod.Data_Mem.F_M.MRAM[26][0] ;
 wire \mod.Data_Mem.F_M.MRAM[26][1] ;
 wire \mod.Data_Mem.F_M.MRAM[26][2] ;
 wire \mod.Data_Mem.F_M.MRAM[26][3] ;
 wire \mod.Data_Mem.F_M.MRAM[26][4] ;
 wire \mod.Data_Mem.F_M.MRAM[26][5] ;
 wire \mod.Data_Mem.F_M.MRAM[26][6] ;
 wire \mod.Data_Mem.F_M.MRAM[26][7] ;
 wire \mod.Data_Mem.F_M.MRAM[27][0] ;
 wire \mod.Data_Mem.F_M.MRAM[27][1] ;
 wire \mod.Data_Mem.F_M.MRAM[27][2] ;
 wire \mod.Data_Mem.F_M.MRAM[27][3] ;
 wire \mod.Data_Mem.F_M.MRAM[27][4] ;
 wire \mod.Data_Mem.F_M.MRAM[27][5] ;
 wire \mod.Data_Mem.F_M.MRAM[27][6] ;
 wire \mod.Data_Mem.F_M.MRAM[27][7] ;
 wire \mod.Data_Mem.F_M.MRAM[28][0] ;
 wire \mod.Data_Mem.F_M.MRAM[28][1] ;
 wire \mod.Data_Mem.F_M.MRAM[28][2] ;
 wire \mod.Data_Mem.F_M.MRAM[28][3] ;
 wire \mod.Data_Mem.F_M.MRAM[28][4] ;
 wire \mod.Data_Mem.F_M.MRAM[28][5] ;
 wire \mod.Data_Mem.F_M.MRAM[28][6] ;
 wire \mod.Data_Mem.F_M.MRAM[28][7] ;
 wire \mod.Data_Mem.F_M.MRAM[29][0] ;
 wire \mod.Data_Mem.F_M.MRAM[29][1] ;
 wire \mod.Data_Mem.F_M.MRAM[29][2] ;
 wire \mod.Data_Mem.F_M.MRAM[29][3] ;
 wire \mod.Data_Mem.F_M.MRAM[29][4] ;
 wire \mod.Data_Mem.F_M.MRAM[29][5] ;
 wire \mod.Data_Mem.F_M.MRAM[29][6] ;
 wire \mod.Data_Mem.F_M.MRAM[29][7] ;
 wire \mod.Data_Mem.F_M.MRAM[2][0] ;
 wire \mod.Data_Mem.F_M.MRAM[2][1] ;
 wire \mod.Data_Mem.F_M.MRAM[2][2] ;
 wire \mod.Data_Mem.F_M.MRAM[2][3] ;
 wire \mod.Data_Mem.F_M.MRAM[2][4] ;
 wire \mod.Data_Mem.F_M.MRAM[2][5] ;
 wire \mod.Data_Mem.F_M.MRAM[2][6] ;
 wire \mod.Data_Mem.F_M.MRAM[2][7] ;
 wire \mod.Data_Mem.F_M.MRAM[30][0] ;
 wire \mod.Data_Mem.F_M.MRAM[30][1] ;
 wire \mod.Data_Mem.F_M.MRAM[30][2] ;
 wire \mod.Data_Mem.F_M.MRAM[30][3] ;
 wire \mod.Data_Mem.F_M.MRAM[30][4] ;
 wire \mod.Data_Mem.F_M.MRAM[30][5] ;
 wire \mod.Data_Mem.F_M.MRAM[30][6] ;
 wire \mod.Data_Mem.F_M.MRAM[30][7] ;
 wire \mod.Data_Mem.F_M.MRAM[31][0] ;
 wire \mod.Data_Mem.F_M.MRAM[31][1] ;
 wire \mod.Data_Mem.F_M.MRAM[31][2] ;
 wire \mod.Data_Mem.F_M.MRAM[31][3] ;
 wire \mod.Data_Mem.F_M.MRAM[31][4] ;
 wire \mod.Data_Mem.F_M.MRAM[31][5] ;
 wire \mod.Data_Mem.F_M.MRAM[31][6] ;
 wire \mod.Data_Mem.F_M.MRAM[31][7] ;
 wire \mod.Data_Mem.F_M.MRAM[3][0] ;
 wire \mod.Data_Mem.F_M.MRAM[3][1] ;
 wire \mod.Data_Mem.F_M.MRAM[3][2] ;
 wire \mod.Data_Mem.F_M.MRAM[3][3] ;
 wire \mod.Data_Mem.F_M.MRAM[3][4] ;
 wire \mod.Data_Mem.F_M.MRAM[3][5] ;
 wire \mod.Data_Mem.F_M.MRAM[3][6] ;
 wire \mod.Data_Mem.F_M.MRAM[3][7] ;
 wire \mod.Data_Mem.F_M.MRAM[4][0] ;
 wire \mod.Data_Mem.F_M.MRAM[4][1] ;
 wire \mod.Data_Mem.F_M.MRAM[4][2] ;
 wire \mod.Data_Mem.F_M.MRAM[4][3] ;
 wire \mod.Data_Mem.F_M.MRAM[4][4] ;
 wire \mod.Data_Mem.F_M.MRAM[4][5] ;
 wire \mod.Data_Mem.F_M.MRAM[4][6] ;
 wire \mod.Data_Mem.F_M.MRAM[4][7] ;
 wire \mod.Data_Mem.F_M.MRAM[5][0] ;
 wire \mod.Data_Mem.F_M.MRAM[5][1] ;
 wire \mod.Data_Mem.F_M.MRAM[5][2] ;
 wire \mod.Data_Mem.F_M.MRAM[5][3] ;
 wire \mod.Data_Mem.F_M.MRAM[5][4] ;
 wire \mod.Data_Mem.F_M.MRAM[5][5] ;
 wire \mod.Data_Mem.F_M.MRAM[5][6] ;
 wire \mod.Data_Mem.F_M.MRAM[5][7] ;
 wire \mod.Data_Mem.F_M.MRAM[6][0] ;
 wire \mod.Data_Mem.F_M.MRAM[6][1] ;
 wire \mod.Data_Mem.F_M.MRAM[6][2] ;
 wire \mod.Data_Mem.F_M.MRAM[6][3] ;
 wire \mod.Data_Mem.F_M.MRAM[6][4] ;
 wire \mod.Data_Mem.F_M.MRAM[6][5] ;
 wire \mod.Data_Mem.F_M.MRAM[6][6] ;
 wire \mod.Data_Mem.F_M.MRAM[6][7] ;
 wire \mod.Data_Mem.F_M.MRAM[768][0] ;
 wire \mod.Data_Mem.F_M.MRAM[768][1] ;
 wire \mod.Data_Mem.F_M.MRAM[768][2] ;
 wire \mod.Data_Mem.F_M.MRAM[768][3] ;
 wire \mod.Data_Mem.F_M.MRAM[768][4] ;
 wire \mod.Data_Mem.F_M.MRAM[768][5] ;
 wire \mod.Data_Mem.F_M.MRAM[768][6] ;
 wire \mod.Data_Mem.F_M.MRAM[768][7] ;
 wire \mod.Data_Mem.F_M.MRAM[769][0] ;
 wire \mod.Data_Mem.F_M.MRAM[769][1] ;
 wire \mod.Data_Mem.F_M.MRAM[769][2] ;
 wire \mod.Data_Mem.F_M.MRAM[769][3] ;
 wire \mod.Data_Mem.F_M.MRAM[769][4] ;
 wire \mod.Data_Mem.F_M.MRAM[769][5] ;
 wire \mod.Data_Mem.F_M.MRAM[769][6] ;
 wire \mod.Data_Mem.F_M.MRAM[769][7] ;
 wire \mod.Data_Mem.F_M.MRAM[770][0] ;
 wire \mod.Data_Mem.F_M.MRAM[770][1] ;
 wire \mod.Data_Mem.F_M.MRAM[770][2] ;
 wire \mod.Data_Mem.F_M.MRAM[770][3] ;
 wire \mod.Data_Mem.F_M.MRAM[770][4] ;
 wire \mod.Data_Mem.F_M.MRAM[770][5] ;
 wire \mod.Data_Mem.F_M.MRAM[770][6] ;
 wire \mod.Data_Mem.F_M.MRAM[770][7] ;
 wire \mod.Data_Mem.F_M.MRAM[771][0] ;
 wire \mod.Data_Mem.F_M.MRAM[771][1] ;
 wire \mod.Data_Mem.F_M.MRAM[771][2] ;
 wire \mod.Data_Mem.F_M.MRAM[771][3] ;
 wire \mod.Data_Mem.F_M.MRAM[771][4] ;
 wire \mod.Data_Mem.F_M.MRAM[771][5] ;
 wire \mod.Data_Mem.F_M.MRAM[771][6] ;
 wire \mod.Data_Mem.F_M.MRAM[771][7] ;
 wire \mod.Data_Mem.F_M.MRAM[772][0] ;
 wire \mod.Data_Mem.F_M.MRAM[772][1] ;
 wire \mod.Data_Mem.F_M.MRAM[772][2] ;
 wire \mod.Data_Mem.F_M.MRAM[772][3] ;
 wire \mod.Data_Mem.F_M.MRAM[772][4] ;
 wire \mod.Data_Mem.F_M.MRAM[772][5] ;
 wire \mod.Data_Mem.F_M.MRAM[772][6] ;
 wire \mod.Data_Mem.F_M.MRAM[772][7] ;
 wire \mod.Data_Mem.F_M.MRAM[773][0] ;
 wire \mod.Data_Mem.F_M.MRAM[773][1] ;
 wire \mod.Data_Mem.F_M.MRAM[773][2] ;
 wire \mod.Data_Mem.F_M.MRAM[773][3] ;
 wire \mod.Data_Mem.F_M.MRAM[773][4] ;
 wire \mod.Data_Mem.F_M.MRAM[773][5] ;
 wire \mod.Data_Mem.F_M.MRAM[773][6] ;
 wire \mod.Data_Mem.F_M.MRAM[773][7] ;
 wire \mod.Data_Mem.F_M.MRAM[774][0] ;
 wire \mod.Data_Mem.F_M.MRAM[774][1] ;
 wire \mod.Data_Mem.F_M.MRAM[774][2] ;
 wire \mod.Data_Mem.F_M.MRAM[774][3] ;
 wire \mod.Data_Mem.F_M.MRAM[774][4] ;
 wire \mod.Data_Mem.F_M.MRAM[774][5] ;
 wire \mod.Data_Mem.F_M.MRAM[774][6] ;
 wire \mod.Data_Mem.F_M.MRAM[774][7] ;
 wire \mod.Data_Mem.F_M.MRAM[775][0] ;
 wire \mod.Data_Mem.F_M.MRAM[775][1] ;
 wire \mod.Data_Mem.F_M.MRAM[775][2] ;
 wire \mod.Data_Mem.F_M.MRAM[775][3] ;
 wire \mod.Data_Mem.F_M.MRAM[775][4] ;
 wire \mod.Data_Mem.F_M.MRAM[775][5] ;
 wire \mod.Data_Mem.F_M.MRAM[775][6] ;
 wire \mod.Data_Mem.F_M.MRAM[775][7] ;
 wire \mod.Data_Mem.F_M.MRAM[776][0] ;
 wire \mod.Data_Mem.F_M.MRAM[776][1] ;
 wire \mod.Data_Mem.F_M.MRAM[776][2] ;
 wire \mod.Data_Mem.F_M.MRAM[776][3] ;
 wire \mod.Data_Mem.F_M.MRAM[776][4] ;
 wire \mod.Data_Mem.F_M.MRAM[776][5] ;
 wire \mod.Data_Mem.F_M.MRAM[776][6] ;
 wire \mod.Data_Mem.F_M.MRAM[776][7] ;
 wire \mod.Data_Mem.F_M.MRAM[777][0] ;
 wire \mod.Data_Mem.F_M.MRAM[777][1] ;
 wire \mod.Data_Mem.F_M.MRAM[777][2] ;
 wire \mod.Data_Mem.F_M.MRAM[777][3] ;
 wire \mod.Data_Mem.F_M.MRAM[777][4] ;
 wire \mod.Data_Mem.F_M.MRAM[777][5] ;
 wire \mod.Data_Mem.F_M.MRAM[777][6] ;
 wire \mod.Data_Mem.F_M.MRAM[777][7] ;
 wire \mod.Data_Mem.F_M.MRAM[778][0] ;
 wire \mod.Data_Mem.F_M.MRAM[778][1] ;
 wire \mod.Data_Mem.F_M.MRAM[778][2] ;
 wire \mod.Data_Mem.F_M.MRAM[778][3] ;
 wire \mod.Data_Mem.F_M.MRAM[778][4] ;
 wire \mod.Data_Mem.F_M.MRAM[778][5] ;
 wire \mod.Data_Mem.F_M.MRAM[778][6] ;
 wire \mod.Data_Mem.F_M.MRAM[778][7] ;
 wire \mod.Data_Mem.F_M.MRAM[779][0] ;
 wire \mod.Data_Mem.F_M.MRAM[779][1] ;
 wire \mod.Data_Mem.F_M.MRAM[779][2] ;
 wire \mod.Data_Mem.F_M.MRAM[779][3] ;
 wire \mod.Data_Mem.F_M.MRAM[779][4] ;
 wire \mod.Data_Mem.F_M.MRAM[779][5] ;
 wire \mod.Data_Mem.F_M.MRAM[779][6] ;
 wire \mod.Data_Mem.F_M.MRAM[779][7] ;
 wire \mod.Data_Mem.F_M.MRAM[780][0] ;
 wire \mod.Data_Mem.F_M.MRAM[780][1] ;
 wire \mod.Data_Mem.F_M.MRAM[780][2] ;
 wire \mod.Data_Mem.F_M.MRAM[780][3] ;
 wire \mod.Data_Mem.F_M.MRAM[780][4] ;
 wire \mod.Data_Mem.F_M.MRAM[780][5] ;
 wire \mod.Data_Mem.F_M.MRAM[780][6] ;
 wire \mod.Data_Mem.F_M.MRAM[780][7] ;
 wire \mod.Data_Mem.F_M.MRAM[781][0] ;
 wire \mod.Data_Mem.F_M.MRAM[781][1] ;
 wire \mod.Data_Mem.F_M.MRAM[781][2] ;
 wire \mod.Data_Mem.F_M.MRAM[781][3] ;
 wire \mod.Data_Mem.F_M.MRAM[781][4] ;
 wire \mod.Data_Mem.F_M.MRAM[781][5] ;
 wire \mod.Data_Mem.F_M.MRAM[781][6] ;
 wire \mod.Data_Mem.F_M.MRAM[781][7] ;
 wire \mod.Data_Mem.F_M.MRAM[782][0] ;
 wire \mod.Data_Mem.F_M.MRAM[782][1] ;
 wire \mod.Data_Mem.F_M.MRAM[782][2] ;
 wire \mod.Data_Mem.F_M.MRAM[782][3] ;
 wire \mod.Data_Mem.F_M.MRAM[782][4] ;
 wire \mod.Data_Mem.F_M.MRAM[782][5] ;
 wire \mod.Data_Mem.F_M.MRAM[782][6] ;
 wire \mod.Data_Mem.F_M.MRAM[782][7] ;
 wire \mod.Data_Mem.F_M.MRAM[783][0] ;
 wire \mod.Data_Mem.F_M.MRAM[783][1] ;
 wire \mod.Data_Mem.F_M.MRAM[783][2] ;
 wire \mod.Data_Mem.F_M.MRAM[783][3] ;
 wire \mod.Data_Mem.F_M.MRAM[783][4] ;
 wire \mod.Data_Mem.F_M.MRAM[783][5] ;
 wire \mod.Data_Mem.F_M.MRAM[783][6] ;
 wire \mod.Data_Mem.F_M.MRAM[783][7] ;
 wire \mod.Data_Mem.F_M.MRAM[784][0] ;
 wire \mod.Data_Mem.F_M.MRAM[784][1] ;
 wire \mod.Data_Mem.F_M.MRAM[784][2] ;
 wire \mod.Data_Mem.F_M.MRAM[784][3] ;
 wire \mod.Data_Mem.F_M.MRAM[784][4] ;
 wire \mod.Data_Mem.F_M.MRAM[784][5] ;
 wire \mod.Data_Mem.F_M.MRAM[784][6] ;
 wire \mod.Data_Mem.F_M.MRAM[784][7] ;
 wire \mod.Data_Mem.F_M.MRAM[785][0] ;
 wire \mod.Data_Mem.F_M.MRAM[785][1] ;
 wire \mod.Data_Mem.F_M.MRAM[785][2] ;
 wire \mod.Data_Mem.F_M.MRAM[785][3] ;
 wire \mod.Data_Mem.F_M.MRAM[785][4] ;
 wire \mod.Data_Mem.F_M.MRAM[785][5] ;
 wire \mod.Data_Mem.F_M.MRAM[785][6] ;
 wire \mod.Data_Mem.F_M.MRAM[785][7] ;
 wire \mod.Data_Mem.F_M.MRAM[786][0] ;
 wire \mod.Data_Mem.F_M.MRAM[786][1] ;
 wire \mod.Data_Mem.F_M.MRAM[786][2] ;
 wire \mod.Data_Mem.F_M.MRAM[786][3] ;
 wire \mod.Data_Mem.F_M.MRAM[786][4] ;
 wire \mod.Data_Mem.F_M.MRAM[786][5] ;
 wire \mod.Data_Mem.F_M.MRAM[786][6] ;
 wire \mod.Data_Mem.F_M.MRAM[786][7] ;
 wire \mod.Data_Mem.F_M.MRAM[787][0] ;
 wire \mod.Data_Mem.F_M.MRAM[787][1] ;
 wire \mod.Data_Mem.F_M.MRAM[787][2] ;
 wire \mod.Data_Mem.F_M.MRAM[787][3] ;
 wire \mod.Data_Mem.F_M.MRAM[787][4] ;
 wire \mod.Data_Mem.F_M.MRAM[787][5] ;
 wire \mod.Data_Mem.F_M.MRAM[787][6] ;
 wire \mod.Data_Mem.F_M.MRAM[787][7] ;
 wire \mod.Data_Mem.F_M.MRAM[788][0] ;
 wire \mod.Data_Mem.F_M.MRAM[788][1] ;
 wire \mod.Data_Mem.F_M.MRAM[788][2] ;
 wire \mod.Data_Mem.F_M.MRAM[788][3] ;
 wire \mod.Data_Mem.F_M.MRAM[788][4] ;
 wire \mod.Data_Mem.F_M.MRAM[788][5] ;
 wire \mod.Data_Mem.F_M.MRAM[788][6] ;
 wire \mod.Data_Mem.F_M.MRAM[788][7] ;
 wire \mod.Data_Mem.F_M.MRAM[789][0] ;
 wire \mod.Data_Mem.F_M.MRAM[789][1] ;
 wire \mod.Data_Mem.F_M.MRAM[789][2] ;
 wire \mod.Data_Mem.F_M.MRAM[789][3] ;
 wire \mod.Data_Mem.F_M.MRAM[789][4] ;
 wire \mod.Data_Mem.F_M.MRAM[789][5] ;
 wire \mod.Data_Mem.F_M.MRAM[789][6] ;
 wire \mod.Data_Mem.F_M.MRAM[789][7] ;
 wire \mod.Data_Mem.F_M.MRAM[790][0] ;
 wire \mod.Data_Mem.F_M.MRAM[790][1] ;
 wire \mod.Data_Mem.F_M.MRAM[790][2] ;
 wire \mod.Data_Mem.F_M.MRAM[790][3] ;
 wire \mod.Data_Mem.F_M.MRAM[790][4] ;
 wire \mod.Data_Mem.F_M.MRAM[790][5] ;
 wire \mod.Data_Mem.F_M.MRAM[790][6] ;
 wire \mod.Data_Mem.F_M.MRAM[790][7] ;
 wire \mod.Data_Mem.F_M.MRAM[791][0] ;
 wire \mod.Data_Mem.F_M.MRAM[791][1] ;
 wire \mod.Data_Mem.F_M.MRAM[791][2] ;
 wire \mod.Data_Mem.F_M.MRAM[791][3] ;
 wire \mod.Data_Mem.F_M.MRAM[791][4] ;
 wire \mod.Data_Mem.F_M.MRAM[791][5] ;
 wire \mod.Data_Mem.F_M.MRAM[791][6] ;
 wire \mod.Data_Mem.F_M.MRAM[791][7] ;
 wire \mod.Data_Mem.F_M.MRAM[792][0] ;
 wire \mod.Data_Mem.F_M.MRAM[792][1] ;
 wire \mod.Data_Mem.F_M.MRAM[792][2] ;
 wire \mod.Data_Mem.F_M.MRAM[792][3] ;
 wire \mod.Data_Mem.F_M.MRAM[792][4] ;
 wire \mod.Data_Mem.F_M.MRAM[792][5] ;
 wire \mod.Data_Mem.F_M.MRAM[792][6] ;
 wire \mod.Data_Mem.F_M.MRAM[792][7] ;
 wire \mod.Data_Mem.F_M.MRAM[793][0] ;
 wire \mod.Data_Mem.F_M.MRAM[793][1] ;
 wire \mod.Data_Mem.F_M.MRAM[793][2] ;
 wire \mod.Data_Mem.F_M.MRAM[793][3] ;
 wire \mod.Data_Mem.F_M.MRAM[793][4] ;
 wire \mod.Data_Mem.F_M.MRAM[793][5] ;
 wire \mod.Data_Mem.F_M.MRAM[793][6] ;
 wire \mod.Data_Mem.F_M.MRAM[793][7] ;
 wire \mod.Data_Mem.F_M.MRAM[794][0] ;
 wire \mod.Data_Mem.F_M.MRAM[794][1] ;
 wire \mod.Data_Mem.F_M.MRAM[794][2] ;
 wire \mod.Data_Mem.F_M.MRAM[794][3] ;
 wire \mod.Data_Mem.F_M.MRAM[794][4] ;
 wire \mod.Data_Mem.F_M.MRAM[794][5] ;
 wire \mod.Data_Mem.F_M.MRAM[794][6] ;
 wire \mod.Data_Mem.F_M.MRAM[794][7] ;
 wire \mod.Data_Mem.F_M.MRAM[795][0] ;
 wire \mod.Data_Mem.F_M.MRAM[795][1] ;
 wire \mod.Data_Mem.F_M.MRAM[795][2] ;
 wire \mod.Data_Mem.F_M.MRAM[795][3] ;
 wire \mod.Data_Mem.F_M.MRAM[795][4] ;
 wire \mod.Data_Mem.F_M.MRAM[795][5] ;
 wire \mod.Data_Mem.F_M.MRAM[795][6] ;
 wire \mod.Data_Mem.F_M.MRAM[795][7] ;
 wire \mod.Data_Mem.F_M.MRAM[796][0] ;
 wire \mod.Data_Mem.F_M.MRAM[796][1] ;
 wire \mod.Data_Mem.F_M.MRAM[796][2] ;
 wire \mod.Data_Mem.F_M.MRAM[796][3] ;
 wire \mod.Data_Mem.F_M.MRAM[796][4] ;
 wire \mod.Data_Mem.F_M.MRAM[796][5] ;
 wire \mod.Data_Mem.F_M.MRAM[796][6] ;
 wire \mod.Data_Mem.F_M.MRAM[796][7] ;
 wire \mod.Data_Mem.F_M.MRAM[797][0] ;
 wire \mod.Data_Mem.F_M.MRAM[797][1] ;
 wire \mod.Data_Mem.F_M.MRAM[797][2] ;
 wire \mod.Data_Mem.F_M.MRAM[797][3] ;
 wire \mod.Data_Mem.F_M.MRAM[797][4] ;
 wire \mod.Data_Mem.F_M.MRAM[797][5] ;
 wire \mod.Data_Mem.F_M.MRAM[797][6] ;
 wire \mod.Data_Mem.F_M.MRAM[797][7] ;
 wire \mod.Data_Mem.F_M.MRAM[798][0] ;
 wire \mod.Data_Mem.F_M.MRAM[798][1] ;
 wire \mod.Data_Mem.F_M.MRAM[798][2] ;
 wire \mod.Data_Mem.F_M.MRAM[798][3] ;
 wire \mod.Data_Mem.F_M.MRAM[798][4] ;
 wire \mod.Data_Mem.F_M.MRAM[798][5] ;
 wire \mod.Data_Mem.F_M.MRAM[798][6] ;
 wire \mod.Data_Mem.F_M.MRAM[798][7] ;
 wire \mod.Data_Mem.F_M.MRAM[799][0] ;
 wire \mod.Data_Mem.F_M.MRAM[799][1] ;
 wire \mod.Data_Mem.F_M.MRAM[799][2] ;
 wire \mod.Data_Mem.F_M.MRAM[799][3] ;
 wire \mod.Data_Mem.F_M.MRAM[799][4] ;
 wire \mod.Data_Mem.F_M.MRAM[799][5] ;
 wire \mod.Data_Mem.F_M.MRAM[799][6] ;
 wire \mod.Data_Mem.F_M.MRAM[799][7] ;
 wire \mod.Data_Mem.F_M.MRAM[7][0] ;
 wire \mod.Data_Mem.F_M.MRAM[7][1] ;
 wire \mod.Data_Mem.F_M.MRAM[7][2] ;
 wire \mod.Data_Mem.F_M.MRAM[7][3] ;
 wire \mod.Data_Mem.F_M.MRAM[7][4] ;
 wire \mod.Data_Mem.F_M.MRAM[7][5] ;
 wire \mod.Data_Mem.F_M.MRAM[7][6] ;
 wire \mod.Data_Mem.F_M.MRAM[7][7] ;
 wire \mod.Data_Mem.F_M.MRAM[8][0] ;
 wire \mod.Data_Mem.F_M.MRAM[8][1] ;
 wire \mod.Data_Mem.F_M.MRAM[8][2] ;
 wire \mod.Data_Mem.F_M.MRAM[8][3] ;
 wire \mod.Data_Mem.F_M.MRAM[8][4] ;
 wire \mod.Data_Mem.F_M.MRAM[8][5] ;
 wire \mod.Data_Mem.F_M.MRAM[8][6] ;
 wire \mod.Data_Mem.F_M.MRAM[8][7] ;
 wire \mod.Data_Mem.F_M.MRAM[9][0] ;
 wire \mod.Data_Mem.F_M.MRAM[9][1] ;
 wire \mod.Data_Mem.F_M.MRAM[9][2] ;
 wire \mod.Data_Mem.F_M.MRAM[9][3] ;
 wire \mod.Data_Mem.F_M.MRAM[9][4] ;
 wire \mod.Data_Mem.F_M.MRAM[9][5] ;
 wire \mod.Data_Mem.F_M.MRAM[9][6] ;
 wire \mod.Data_Mem.F_M.MRAM[9][7] ;
 wire \mod.Data_Mem.F_M.dest[0] ;
 wire \mod.Data_Mem.F_M.dest[1] ;
 wire \mod.Data_Mem.F_M.dest[2] ;
 wire \mod.Data_Mem.F_M.dest[4] ;
 wire \mod.Data_Mem.F_M.dest[8] ;
 wire \mod.Data_Mem.F_M.out_data[0] ;
 wire \mod.Data_Mem.F_M.out_data[10] ;
 wire \mod.Data_Mem.F_M.out_data[11] ;
 wire \mod.Data_Mem.F_M.out_data[12] ;
 wire \mod.Data_Mem.F_M.out_data[13] ;
 wire \mod.Data_Mem.F_M.out_data[14] ;
 wire \mod.Data_Mem.F_M.out_data[15] ;
 wire \mod.Data_Mem.F_M.out_data[16] ;
 wire \mod.Data_Mem.F_M.out_data[17] ;
 wire \mod.Data_Mem.F_M.out_data[18] ;
 wire \mod.Data_Mem.F_M.out_data[19] ;
 wire \mod.Data_Mem.F_M.out_data[1] ;
 wire \mod.Data_Mem.F_M.out_data[20] ;
 wire \mod.Data_Mem.F_M.out_data[21] ;
 wire \mod.Data_Mem.F_M.out_data[22] ;
 wire \mod.Data_Mem.F_M.out_data[23] ;
 wire \mod.Data_Mem.F_M.out_data[24] ;
 wire \mod.Data_Mem.F_M.out_data[25] ;
 wire \mod.Data_Mem.F_M.out_data[26] ;
 wire \mod.Data_Mem.F_M.out_data[27] ;
 wire \mod.Data_Mem.F_M.out_data[28] ;
 wire \mod.Data_Mem.F_M.out_data[29] ;
 wire \mod.Data_Mem.F_M.out_data[2] ;
 wire \mod.Data_Mem.F_M.out_data[30] ;
 wire \mod.Data_Mem.F_M.out_data[31] ;
 wire \mod.Data_Mem.F_M.out_data[32] ;
 wire \mod.Data_Mem.F_M.out_data[33] ;
 wire \mod.Data_Mem.F_M.out_data[34] ;
 wire \mod.Data_Mem.F_M.out_data[35] ;
 wire \mod.Data_Mem.F_M.out_data[36] ;
 wire \mod.Data_Mem.F_M.out_data[37] ;
 wire \mod.Data_Mem.F_M.out_data[38] ;
 wire \mod.Data_Mem.F_M.out_data[39] ;
 wire \mod.Data_Mem.F_M.out_data[3] ;
 wire \mod.Data_Mem.F_M.out_data[40] ;
 wire \mod.Data_Mem.F_M.out_data[41] ;
 wire \mod.Data_Mem.F_M.out_data[42] ;
 wire \mod.Data_Mem.F_M.out_data[43] ;
 wire \mod.Data_Mem.F_M.out_data[44] ;
 wire \mod.Data_Mem.F_M.out_data[45] ;
 wire \mod.Data_Mem.F_M.out_data[46] ;
 wire \mod.Data_Mem.F_M.out_data[47] ;
 wire \mod.Data_Mem.F_M.out_data[48] ;
 wire \mod.Data_Mem.F_M.out_data[49] ;
 wire \mod.Data_Mem.F_M.out_data[4] ;
 wire \mod.Data_Mem.F_M.out_data[50] ;
 wire \mod.Data_Mem.F_M.out_data[51] ;
 wire \mod.Data_Mem.F_M.out_data[52] ;
 wire \mod.Data_Mem.F_M.out_data[53] ;
 wire \mod.Data_Mem.F_M.out_data[54] ;
 wire \mod.Data_Mem.F_M.out_data[55] ;
 wire \mod.Data_Mem.F_M.out_data[56] ;
 wire \mod.Data_Mem.F_M.out_data[57] ;
 wire \mod.Data_Mem.F_M.out_data[58] ;
 wire \mod.Data_Mem.F_M.out_data[59] ;
 wire \mod.Data_Mem.F_M.out_data[5] ;
 wire \mod.Data_Mem.F_M.out_data[60] ;
 wire \mod.Data_Mem.F_M.out_data[61] ;
 wire \mod.Data_Mem.F_M.out_data[62] ;
 wire \mod.Data_Mem.F_M.out_data[63] ;
 wire \mod.Data_Mem.F_M.out_data[64] ;
 wire \mod.Data_Mem.F_M.out_data[65] ;
 wire \mod.Data_Mem.F_M.out_data[66] ;
 wire \mod.Data_Mem.F_M.out_data[67] ;
 wire \mod.Data_Mem.F_M.out_data[68] ;
 wire \mod.Data_Mem.F_M.out_data[69] ;
 wire \mod.Data_Mem.F_M.out_data[6] ;
 wire \mod.Data_Mem.F_M.out_data[70] ;
 wire \mod.Data_Mem.F_M.out_data[71] ;
 wire \mod.Data_Mem.F_M.out_data[72] ;
 wire \mod.Data_Mem.F_M.out_data[73] ;
 wire \mod.Data_Mem.F_M.out_data[74] ;
 wire \mod.Data_Mem.F_M.out_data[75] ;
 wire \mod.Data_Mem.F_M.out_data[76] ;
 wire \mod.Data_Mem.F_M.out_data[77] ;
 wire \mod.Data_Mem.F_M.out_data[78] ;
 wire \mod.Data_Mem.F_M.out_data[79] ;
 wire \mod.Data_Mem.F_M.out_data[7] ;
 wire \mod.Data_Mem.F_M.out_data[8] ;
 wire \mod.Data_Mem.F_M.out_data[9] ;
 wire \mod.Data_Mem.F_M.src[0] ;
 wire \mod.Data_Mem.F_M.src[1] ;
 wire \mod.Data_Mem.F_M.src[2] ;
 wire \mod.Data_Mem.F_M.src[4] ;
 wire \mod.Data_Mem.F_M.src[8] ;
 wire \mod.I_addr[0] ;
 wire \mod.I_addr[1] ;
 wire \mod.I_addr[2] ;
 wire \mod.I_addr[3] ;
 wire \mod.I_addr[4] ;
 wire \mod.I_addr[5] ;
 wire \mod.I_addr[6] ;
 wire \mod.I_addr[7] ;
 wire \mod.Instr_Mem.instruction[10] ;
 wire \mod.Instr_Mem.instruction[11] ;
 wire \mod.Instr_Mem.instruction[13] ;
 wire \mod.Instr_Mem.instruction[17] ;
 wire \mod.Instr_Mem.instruction[22] ;
 wire \mod.Instr_Mem.instruction[23] ;
 wire \mod.Instr_Mem.instruction[24] ;
 wire \mod.Instr_Mem.instruction[26] ;
 wire \mod.Instr_Mem.instruction[30] ;
 wire \mod.Instr_Mem.instruction[7] ;
 wire \mod.Instr_Mem.instruction[8] ;
 wire \mod.Instr_Mem.instruction[9] ;
 wire \mod.P1.instr_reg[10] ;
 wire \mod.P1.instr_reg[11] ;
 wire \mod.P1.instr_reg[13] ;
 wire \mod.P1.instr_reg[17] ;
 wire \mod.P1.instr_reg[7] ;
 wire \mod.P1.instr_reg[8] ;
 wire \mod.P1.instr_reg[9] ;
 wire \mod.P2.Rout_reg1[0] ;
 wire \mod.P2.Rout_reg1[1] ;
 wire \mod.P2.Rout_reg[0] ;
 wire \mod.P2.Rout_reg[1] ;
 wire \mod.P2.dest_reg1[0] ;
 wire \mod.P2.dest_reg1[1] ;
 wire \mod.P2.dest_reg1[2] ;
 wire \mod.P2.dest_reg1[4] ;
 wire \mod.P2.dest_reg1[8] ;
 wire \mod.P2.dest_reg[0] ;
 wire \mod.P2.dest_reg[1] ;
 wire \mod.P2.dest_reg[2] ;
 wire \mod.P2.dest_reg[4] ;
 wire \mod.P2.dest_reg[8] ;
 wire \mod.P3.Res[0] ;
 wire \mod.P3.Res[1] ;
 wire \mod.P3.Res[2] ;
 wire \mod.P3.Res[3] ;
 wire \mod.P3.Res[4] ;
 wire \mod.P3.Res[5] ;
 wire \mod.P3.Res[6] ;
 wire \mod.P3.Res[7] ;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net149;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net150;
 wire net178;
 wire net179;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;

 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3933_ (.I(\mod.I_addr[0] ),
    .Z(_0612_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3934_ (.I(_0612_),
    .ZN(_0080_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3935_ (.I(\mod.Arithmetic.CN.F_in[0] ),
    .Z(_0613_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3936_ (.I(_0613_),
    .Z(_0614_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3937_ (.I(_0614_),
    .Z(_0615_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3938_ (.I(_0615_),
    .Z(_0616_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3939_ (.I(_0616_),
    .Z(_0617_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3940_ (.I(_0617_),
    .Z(_0618_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3941_ (.I(_0618_),
    .Z(_0619_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3942_ (.I(_0619_),
    .Z(_0620_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3943_ (.I(_0620_),
    .Z(_0621_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3944_ (.I(_0621_),
    .Z(_0622_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3945_ (.I(_0622_),
    .Z(_0623_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3946_ (.I(_0623_),
    .Z(_0624_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3947_ (.I(_0624_),
    .Z(_0625_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _3948_ (.A1(\mod.P1.instr_reg[17] ),
    .A2(_0625_),
    .Z(_0626_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3949_ (.I(_0626_),
    .Z(\mod.DM_en ));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3950_ (.A1(\mod.P2.Rout_reg[0] ),
    .A2(\mod.P2.Rout_reg[1] ),
    .ZN(_0627_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3951_ (.I(_0627_),
    .Z(_0628_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3952_ (.I(_0628_),
    .Z(_0629_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3953_ (.I(\mod.Arithmetic.CN.I_in[8] ),
    .Z(_0630_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3954_ (.A1(_0622_),
    .A2(_0630_),
    .ZN(_0631_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3955_ (.I(_0613_),
    .Z(_0632_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3956_ (.I(_0632_),
    .Z(_0633_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _3957_ (.I(_0633_),
    .Z(_0634_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3958_ (.I(_0634_),
    .Z(_0635_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3959_ (.I(_0635_),
    .Z(_0636_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3960_ (.I(_0636_),
    .Z(_0637_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3961_ (.I(\mod.Arithmetic.CN.I_in[16] ),
    .Z(_0638_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _3962_ (.A1(_0637_),
    .A2(\mod.Arithmetic.CN.I_in[24] ),
    .A3(_0638_),
    .ZN(_0639_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3963_ (.I(_0613_),
    .Z(_0640_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3964_ (.I(_0640_),
    .Z(_0641_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3965_ (.I(_0641_),
    .Z(_0642_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3966_ (.I(_0642_),
    .Z(_0643_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3967_ (.A1(_0643_),
    .A2(\mod.Arithmetic.CN.I_in[16] ),
    .ZN(_0644_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3968_ (.I(_0641_),
    .Z(_0645_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3969_ (.A1(_0645_),
    .A2(\mod.Arithmetic.CN.I_in[24] ),
    .ZN(_0646_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3970_ (.A1(_0644_),
    .A2(_0646_),
    .ZN(_0647_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3971_ (.A1(_0639_),
    .A2(_0647_),
    .ZN(_0648_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _3972_ (.A1(_0631_),
    .A2(_0648_),
    .Z(_0649_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3973_ (.I(_0645_),
    .Z(_0650_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3974_ (.I(_0650_),
    .Z(_0651_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3975_ (.A1(_0651_),
    .A2(\mod.Arithmetic.CN.I_in[32] ),
    .ZN(_0652_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3976_ (.I(_0616_),
    .Z(_0653_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3977_ (.I(_0653_),
    .Z(_0654_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3978_ (.I(_0654_),
    .Z(_0655_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3979_ (.I(\mod.Arithmetic.CN.I_in[40] ),
    .Z(_0656_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3980_ (.A1(_0655_),
    .A2(_0656_),
    .ZN(_0657_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _3981_ (.A1(_0636_),
    .A2(\mod.Arithmetic.CN.I_in[48] ),
    .ZN(_0658_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3982_ (.A1(_0635_),
    .A2(\mod.Arithmetic.CN.I_in[56] ),
    .ZN(_0659_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3983_ (.I(_0659_),
    .Z(_0660_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3984_ (.I(\mod.Arithmetic.ACTI.x[0] ),
    .Z(_0661_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _3985_ (.A1(_0650_),
    .A2(_0661_),
    .A3(\mod.Arithmetic.CN.I_in[64] ),
    .ZN(_0662_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3986_ (.A1(_0640_),
    .A2(\mod.Arithmetic.CN.I_in[64] ),
    .ZN(_0663_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3987_ (.A1(_0633_),
    .A2(\mod.Arithmetic.ACTI.x[0] ),
    .ZN(_0664_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3988_ (.I(_0664_),
    .Z(_0665_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3989_ (.A1(_0663_),
    .A2(_0665_),
    .ZN(_0666_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3990_ (.A1(_0662_),
    .A2(_0666_),
    .ZN(_0667_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _3991_ (.A1(_0660_),
    .A2(_0667_),
    .Z(_0668_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _3992_ (.A1(_0658_),
    .A2(_0668_),
    .ZN(_0669_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _3993_ (.A1(_0652_),
    .A2(_0657_),
    .A3(_0669_),
    .Z(_0670_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _3994_ (.A1(_0649_),
    .A2(_0670_),
    .ZN(_0671_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3995_ (.I(\mod.P2.Rout_reg[1] ),
    .Z(_0672_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _3996_ (.I(\mod.Arithmetic.ACTI.x[7] ),
    .Z(_0673_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3997_ (.I(\mod.Arithmetic.CN.I_in[23] ),
    .Z(_0674_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3998_ (.I(\mod.Arithmetic.CN.I_in[15] ),
    .Z(_0675_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _3999_ (.A1(_0674_),
    .A2(\mod.Arithmetic.I_out[79] ),
    .A3(_0675_),
    .ZN(_0676_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _4000_ (.I(\mod.Arithmetic.I_out[79] ),
    .ZN(_0677_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4001_ (.I(\mod.Arithmetic.CN.I_in[21] ),
    .Z(_0678_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _4002_ (.I(_0678_),
    .ZN(_0679_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _4003_ (.I(\mod.Arithmetic.CN.I_in[19] ),
    .Z(_0680_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _4004_ (.I(\mod.Arithmetic.I_out[75] ),
    .ZN(_0681_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4005_ (.I(\mod.Arithmetic.CN.I_in[18] ),
    .Z(_0682_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _4006_ (.I(\mod.Arithmetic.I_out[74] ),
    .ZN(_0683_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _4007_ (.I(\mod.Arithmetic.CN.I_in[17] ),
    .ZN(_0684_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _4008_ (.I(_0638_),
    .ZN(_0685_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_4 _4009_ (.A1(_0684_),
    .A2(\mod.Arithmetic.I_out[73] ),
    .B(\mod.Arithmetic.I_out[72] ),
    .C(_0685_),
    .ZN(_0686_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _4010_ (.I(_0682_),
    .ZN(_0687_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_2 _4011_ (.A1(_0687_),
    .A2(\mod.Arithmetic.I_out[74] ),
    .B1(_0684_),
    .B2(\mod.Arithmetic.I_out[73] ),
    .ZN(_0688_));
 gf180mcu_fd_sc_mcu7t5v0__oai222_4 _4012_ (.A1(_0680_),
    .A2(_0681_),
    .B1(_0682_),
    .B2(_0683_),
    .C1(_0686_),
    .C2(_0688_),
    .ZN(_0689_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4013_ (.I(\mod.Arithmetic.I_out[76] ),
    .ZN(_0690_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4014_ (.I(\mod.Arithmetic.CN.I_in[20] ),
    .Z(_0691_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _4015_ (.A1(_0690_),
    .A2(_0691_),
    .B1(_0680_),
    .B2(_0681_),
    .ZN(_0692_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4016_ (.A1(_0690_),
    .A2(_0691_),
    .ZN(_0693_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _4017_ (.A1(_0679_),
    .A2(\mod.Arithmetic.I_out[77] ),
    .B1(_0689_),
    .B2(_0692_),
    .C(_0693_),
    .ZN(_0694_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4018_ (.I(\mod.Arithmetic.CN.I_in[22] ),
    .ZN(_0695_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _4019_ (.I(_0695_),
    .Z(_0696_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _4020_ (.A1(\mod.Arithmetic.CN.I_in[23] ),
    .A2(_0677_),
    .ZN(_0697_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4021_ (.I(\mod.Arithmetic.I_out[77] ),
    .ZN(_0698_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _4022_ (.A1(_0696_),
    .A2(\mod.Arithmetic.I_out[78] ),
    .B1(_0678_),
    .B2(_0698_),
    .ZN(_0699_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_4 _4023_ (.A1(_0696_),
    .A2(\mod.Arithmetic.I_out[78] ),
    .B(_0697_),
    .C(_0699_),
    .ZN(_0700_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _4024_ (.A1(_0696_),
    .A2(\mod.Arithmetic.I_out[78] ),
    .A3(_0697_),
    .ZN(_0701_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_4 _4025_ (.A1(\mod.Arithmetic.CN.I_in[23] ),
    .A2(_0677_),
    .B1(_0694_),
    .B2(_0700_),
    .C(_0701_),
    .ZN(_0702_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _4026_ (.I(_0702_),
    .Z(_0703_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _4027_ (.I0(_0638_),
    .I1(\mod.Arithmetic.I_out[72] ),
    .S(_0703_),
    .Z(_0704_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4028_ (.A1(_0674_),
    .A2(\mod.Arithmetic.I_out[79] ),
    .ZN(_0705_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _4029_ (.A1(_0675_),
    .A2(_0705_),
    .Z(_0706_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4030_ (.I(\mod.Arithmetic.CN.I_in[10] ),
    .ZN(_0707_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _4031_ (.I0(_0682_),
    .I1(\mod.Arithmetic.I_out[74] ),
    .S(_0703_),
    .Z(_0708_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4032_ (.I(\mod.Arithmetic.CN.I_in[9] ),
    .Z(_0709_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4033_ (.I(_0709_),
    .Z(_0710_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4034_ (.I(\mod.Arithmetic.I_out[73] ),
    .ZN(_0711_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _4035_ (.I0(_0684_),
    .I1(_0711_),
    .S(_0702_),
    .Z(_0712_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _4036_ (.I(_0702_),
    .Z(_0713_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _4037_ (.I0(_0687_),
    .I1(_0683_),
    .S(_0713_),
    .Z(_0714_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4038_ (.I(\mod.Arithmetic.CN.I_in[10] ),
    .Z(_0715_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4039_ (.I(_0715_),
    .Z(_0716_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4040_ (.A1(_0710_),
    .A2(_0712_),
    .B1(_0714_),
    .B2(_0716_),
    .ZN(_0717_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4041_ (.I(\mod.Arithmetic.I_out[72] ),
    .ZN(_0718_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _4042_ (.I0(_0685_),
    .I1(_0718_),
    .S(_0702_),
    .Z(_0719_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4043_ (.A1(_0710_),
    .A2(_0712_),
    .B(_0719_),
    .C(_0630_),
    .ZN(_0720_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _4044_ (.I0(_0680_),
    .I1(\mod.Arithmetic.I_out[75] ),
    .S(_0713_),
    .Z(_0721_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _4045_ (.I(\mod.Arithmetic.CN.I_in[11] ),
    .ZN(_0722_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _4046_ (.A1(_0707_),
    .A2(_0708_),
    .B1(_0717_),
    .B2(_0720_),
    .C1(_0721_),
    .C2(_0722_),
    .ZN(_0723_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4047_ (.I(\mod.Arithmetic.CN.I_in[12] ),
    .Z(_0724_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4048_ (.I(_0724_),
    .Z(_0725_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4049_ (.I(_0691_),
    .ZN(_0726_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _4050_ (.I0(_0726_),
    .I1(_0690_),
    .S(_0713_),
    .Z(_0727_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _4051_ (.A1(_0725_),
    .A2(_0727_),
    .Z(_0728_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4052_ (.A1(_0722_),
    .A2(_0721_),
    .ZN(_0729_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _4053_ (.I0(_0679_),
    .I1(_0698_),
    .S(_0713_),
    .Z(_0730_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4054_ (.I(\mod.Arithmetic.CN.I_in[13] ),
    .Z(_0731_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _4055_ (.A1(_0725_),
    .A2(_0727_),
    .B1(_0730_),
    .B2(_0731_),
    .ZN(_0732_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4056_ (.I(_0732_),
    .ZN(_0733_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _4057_ (.A1(_0723_),
    .A2(_0728_),
    .A3(_0729_),
    .B(_0733_),
    .ZN(_0734_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4058_ (.I(_0731_),
    .Z(_0735_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4059_ (.A1(_0735_),
    .A2(_0730_),
    .ZN(_0736_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4060_ (.I(\mod.Arithmetic.CN.I_in[14] ),
    .Z(_0737_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _4061_ (.A1(_0674_),
    .A2(_0677_),
    .B1(_0694_),
    .B2(_0700_),
    .ZN(_0738_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4062_ (.I(_0738_),
    .ZN(_0739_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_2 _4063_ (.A1(\mod.Arithmetic.I_out[78] ),
    .A2(_0739_),
    .B1(_0703_),
    .B2(\mod.Arithmetic.CN.I_in[22] ),
    .ZN(_0740_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4064_ (.A1(_0737_),
    .A2(_0740_),
    .ZN(_0741_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _4065_ (.A1(_0736_),
    .A2(_0741_),
    .Z(_0742_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4066_ (.I(_0737_),
    .Z(_0743_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _4067_ (.A1(\mod.Arithmetic.CN.I_in[15] ),
    .A2(_0705_),
    .B1(_0740_),
    .B2(_0743_),
    .ZN(_0744_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _4068_ (.A1(_0734_),
    .A2(_0742_),
    .B(_0744_),
    .ZN(_0745_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _4069_ (.A1(_0706_),
    .A2(_0745_),
    .ZN(_0746_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _4070_ (.I0(_0630_),
    .I1(_0704_),
    .S(_0746_),
    .Z(_0747_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4071_ (.I(\mod.Arithmetic.ACTI.x[1] ),
    .Z(_0748_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4072_ (.A1(_0675_),
    .A2(_0705_),
    .ZN(_0749_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4073_ (.I(_0710_),
    .ZN(_0750_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _4074_ (.I0(\mod.Arithmetic.CN.I_in[17] ),
    .I1(\mod.Arithmetic.I_out[73] ),
    .S(_0703_),
    .Z(_0751_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4075_ (.I(_0630_),
    .ZN(_0752_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _4076_ (.A1(_0750_),
    .A2(_0751_),
    .B(_0704_),
    .C(_0752_),
    .ZN(_0753_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4077_ (.I(_0707_),
    .Z(_0754_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _4078_ (.A1(_0750_),
    .A2(_0751_),
    .B1(_0708_),
    .B2(_0754_),
    .ZN(_0755_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4079_ (.A1(_0754_),
    .A2(_0708_),
    .B1(_0721_),
    .B2(_0722_),
    .ZN(_0756_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4080_ (.A1(_0753_),
    .A2(_0755_),
    .B(_0756_),
    .ZN(_0757_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4081_ (.A1(_0728_),
    .A2(_0729_),
    .ZN(_0758_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4082_ (.A1(_0757_),
    .A2(_0758_),
    .B(_0732_),
    .ZN(_0759_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4083_ (.A1(_0736_),
    .A2(_0741_),
    .ZN(_0760_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4084_ (.I(_0744_),
    .ZN(_0761_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4085_ (.A1(_0759_),
    .A2(_0760_),
    .B(_0761_),
    .ZN(_0762_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4086_ (.A1(_0749_),
    .A2(_0762_),
    .B(_0710_),
    .ZN(_0763_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _4087_ (.A1(_0706_),
    .A2(_0751_),
    .A3(_0745_),
    .ZN(_0764_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _4088_ (.A1(_0748_),
    .A2(_0763_),
    .A3(_0764_),
    .B(_0661_),
    .ZN(_0765_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4089_ (.I(_0746_),
    .Z(_0766_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _4090_ (.A1(_0749_),
    .A2(_0708_),
    .A3(_0762_),
    .ZN(_0767_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4091_ (.I(\mod.Arithmetic.ACTI.x[2] ),
    .Z(_0768_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4092_ (.A1(_0754_),
    .A2(_0766_),
    .B(_0767_),
    .C(_0768_),
    .ZN(_0769_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4093_ (.A1(_0763_),
    .A2(_0764_),
    .B(_0748_),
    .ZN(_0770_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4094_ (.A1(_0747_),
    .A2(_0765_),
    .B(_0769_),
    .C(_0770_),
    .ZN(_0771_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4095_ (.I(_0768_),
    .ZN(_0772_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4096_ (.A1(_0754_),
    .A2(_0766_),
    .B(_0767_),
    .ZN(_0773_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _4097_ (.I0(\mod.Arithmetic.CN.I_in[11] ),
    .I1(_0721_),
    .S(_0746_),
    .Z(_0774_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4098_ (.I(\mod.Arithmetic.ACTI.x[3] ),
    .Z(_0775_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4099_ (.I(_0775_),
    .ZN(_0776_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4100_ (.A1(_0772_),
    .A2(_0773_),
    .B1(_0774_),
    .B2(_0776_),
    .ZN(_0777_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4101_ (.I(_0746_),
    .Z(_0778_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4102_ (.A1(_0727_),
    .A2(_0766_),
    .ZN(_0779_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _4103_ (.A1(_0725_),
    .A2(_0778_),
    .B(_0779_),
    .ZN(_0780_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4104_ (.I(\mod.Arithmetic.ACTI.x[4] ),
    .Z(_0781_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4105_ (.A1(_0776_),
    .A2(_0774_),
    .ZN(_0782_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _4106_ (.A1(_0771_),
    .A2(_0777_),
    .B1(_0780_),
    .B2(_0781_),
    .C(_0782_),
    .ZN(_0783_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4107_ (.A1(_0730_),
    .A2(_0778_),
    .ZN(_0784_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4108_ (.A1(_0735_),
    .A2(_0778_),
    .B(_0784_),
    .ZN(_0785_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4109_ (.I(\mod.Arithmetic.ACTI.x[5] ),
    .Z(_0786_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _4110_ (.A1(_0781_),
    .A2(_0780_),
    .B1(_0785_),
    .B2(_0786_),
    .ZN(_0787_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4111_ (.A1(_0740_),
    .A2(_0766_),
    .ZN(_0788_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4112_ (.A1(_0743_),
    .A2(_0778_),
    .B(_0788_),
    .ZN(_0789_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4113_ (.A1(_0786_),
    .A2(_0785_),
    .B1(_0789_),
    .B2(\mod.Arithmetic.ACTI.x[6] ),
    .ZN(_0790_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _4114_ (.A1(_0783_),
    .A2(_0787_),
    .B(_0790_),
    .ZN(_0791_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _4115_ (.A1(\mod.Arithmetic.ACTI.x[7] ),
    .A2(_0676_),
    .B1(_0789_),
    .B2(\mod.Arithmetic.ACTI.x[6] ),
    .ZN(_0792_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4116_ (.I(_0792_),
    .ZN(_0793_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _4117_ (.A1(_0673_),
    .A2(_0676_),
    .B1(_0791_),
    .B2(_0793_),
    .ZN(_0794_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4118_ (.I(_0794_),
    .Z(_0795_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _4119_ (.A1(_0672_),
    .A2(_0673_),
    .B1(_0795_),
    .B2(\mod.P2.Rout_reg[0] ),
    .ZN(_0796_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4120_ (.I(\mod.P2.Rout_reg[0] ),
    .ZN(_0797_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _4121_ (.A1(_0797_),
    .A2(_0747_),
    .Z(_0798_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4122_ (.I(_0794_),
    .Z(_0799_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _4123_ (.A1(_0661_),
    .A2(_0796_),
    .B1(_0798_),
    .B2(_0799_),
    .C(_0628_),
    .ZN(_0800_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4124_ (.A1(_0629_),
    .A2(_0671_),
    .B(_0800_),
    .ZN(\mod.P3.Res[0] ));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _4125_ (.A1(_0649_),
    .A2(_0670_),
    .Z(_0801_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4126_ (.A1(_0631_),
    .A2(_0648_),
    .ZN(_0802_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4127_ (.A1(_0633_),
    .A2(\mod.Arithmetic.CN.I_in[17] ),
    .ZN(_0803_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4128_ (.I(_0803_),
    .Z(_0804_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4129_ (.I(_0804_),
    .ZN(_0805_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4130_ (.I(\mod.Arithmetic.CN.F_in[0] ),
    .Z(_0806_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4131_ (.I(_0806_),
    .Z(_0807_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4132_ (.A1(_0807_),
    .A2(\mod.Arithmetic.CN.I_in[25] ),
    .ZN(_0808_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4133_ (.I(_0808_),
    .Z(_0809_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4134_ (.A1(_0646_),
    .A2(_0809_),
    .Z(_0810_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _4135_ (.A1(_0644_),
    .A2(_0805_),
    .A3(_0810_),
    .Z(_0811_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _4136_ (.A1(_0639_),
    .A2(_0811_),
    .ZN(_0812_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4137_ (.I(_0637_),
    .Z(_0813_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4138_ (.A1(_0813_),
    .A2(_0709_),
    .ZN(_0814_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4139_ (.A1(_0631_),
    .A2(_0814_),
    .ZN(_0815_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _4140_ (.A1(_0621_),
    .A2(\mod.Arithmetic.CN.I_in[8] ),
    .A3(_0709_),
    .ZN(_0816_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4141_ (.A1(_0815_),
    .A2(_0816_),
    .ZN(_0817_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4142_ (.A1(_0812_),
    .A2(_0817_),
    .Z(_0818_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4143_ (.A1(_0802_),
    .A2(_0818_),
    .Z(_0819_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4144_ (.I(\mod.Arithmetic.CN.I_in[32] ),
    .Z(_0820_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _4145_ (.A1(_0621_),
    .A2(_0656_),
    .A3(_0820_),
    .ZN(_0821_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4146_ (.A1(_0652_),
    .A2(_0657_),
    .ZN(_0822_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _4147_ (.A1(_0821_),
    .A2(_0822_),
    .A3(_0669_),
    .ZN(_0823_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4148_ (.I(_0620_),
    .Z(_0824_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _4149_ (.A1(_0824_),
    .A2(\mod.Arithmetic.CN.I_in[48] ),
    .A3(_0668_),
    .ZN(_0825_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _4150_ (.A1(_0651_),
    .A2(\mod.Arithmetic.CN.I_in[33] ),
    .ZN(_0826_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4151_ (.A1(_0652_),
    .A2(_0826_),
    .ZN(_0827_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _4152_ (.I(_0618_),
    .Z(_0828_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _4153_ (.A1(_0828_),
    .A2(_0820_),
    .A3(\mod.Arithmetic.CN.I_in[33] ),
    .ZN(_0829_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4154_ (.A1(_0827_),
    .A2(_0829_),
    .ZN(_0830_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4155_ (.A1(_0655_),
    .A2(\mod.Arithmetic.CN.I_in[41] ),
    .ZN(_0831_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4156_ (.A1(_0657_),
    .A2(_0831_),
    .ZN(_0832_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _4157_ (.A1(_0655_),
    .A2(\mod.Arithmetic.CN.I_in[40] ),
    .A3(\mod.Arithmetic.CN.I_in[41] ),
    .ZN(_0833_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4158_ (.A1(_0832_),
    .A2(_0833_),
    .ZN(_0834_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4159_ (.A1(_0830_),
    .A2(_0834_),
    .Z(_0835_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _4160_ (.A1(_0821_),
    .A2(_0835_),
    .ZN(_0836_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4161_ (.A1(_0660_),
    .A2(_0667_),
    .ZN(_0837_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4162_ (.A1(_0635_),
    .A2(\mod.Arithmetic.CN.I_in[49] ),
    .ZN(_0838_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _4163_ (.A1(_0658_),
    .A2(_0838_),
    .ZN(_0839_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4164_ (.A1(_0617_),
    .A2(\mod.Arithmetic.CN.I_in[57] ),
    .ZN(_0840_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _4165_ (.A1(_0659_),
    .A2(_0840_),
    .ZN(_0841_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4166_ (.A1(_0807_),
    .A2(\mod.Arithmetic.CN.I_in[65] ),
    .ZN(_0842_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4167_ (.I(\mod.Arithmetic.CN.F_in[0] ),
    .Z(_0843_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4168_ (.I(_0843_),
    .Z(_0844_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4169_ (.A1(_0844_),
    .A2(\mod.Arithmetic.ACTI.x[1] ),
    .ZN(_0845_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _4170_ (.A1(_0663_),
    .A2(_0845_),
    .ZN(_0846_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _4171_ (.A1(_0665_),
    .A2(_0842_),
    .A3(_0846_),
    .ZN(_0847_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _4172_ (.A1(_0662_),
    .A2(_0841_),
    .A3(_0847_),
    .Z(_0848_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _4173_ (.A1(_0837_),
    .A2(_0839_),
    .A3(_0848_),
    .Z(_0849_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _4174_ (.A1(_0825_),
    .A2(_0836_),
    .A3(_0849_),
    .Z(_0850_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _4175_ (.A1(_0823_),
    .A2(_0850_),
    .ZN(_0851_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4176_ (.A1(_0819_),
    .A2(_0851_),
    .Z(_0852_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _4177_ (.A1(_0801_),
    .A2(_0852_),
    .ZN(_0853_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4178_ (.A1(_0672_),
    .A2(_0673_),
    .ZN(_0854_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4179_ (.I(_0854_),
    .Z(_0855_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _4180_ (.A1(_0797_),
    .A2(\mod.P2.Rout_reg[1] ),
    .Z(_0856_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4181_ (.I(_0856_),
    .Z(_0857_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4182_ (.A1(_0763_),
    .A2(_0764_),
    .ZN(_0858_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _4183_ (.I0(_0748_),
    .I1(_0858_),
    .S(_0795_),
    .Z(_0859_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _4184_ (.A1(_0748_),
    .A2(_0855_),
    .B1(_0857_),
    .B2(_0859_),
    .C(_0628_),
    .ZN(_0860_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4185_ (.A1(_0629_),
    .A2(_0853_),
    .B(_0860_),
    .ZN(\mod.P3.Res[1] ));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4186_ (.A1(_0801_),
    .A2(_0852_),
    .ZN(_0861_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4187_ (.A1(_0802_),
    .A2(_0818_),
    .ZN(_0862_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _4188_ (.A1(_0821_),
    .A2(_0822_),
    .A3(_0669_),
    .A4(_0850_),
    .ZN(_0863_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4189_ (.A1(_0819_),
    .A2(_0851_),
    .ZN(_0864_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4190_ (.A1(_0863_),
    .A2(_0864_),
    .ZN(_0865_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4191_ (.A1(_0812_),
    .A2(_0817_),
    .ZN(_0866_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _4192_ (.A1(_0623_),
    .A2(_0656_),
    .A3(_0820_),
    .A4(_0835_),
    .ZN(_0867_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4193_ (.A1(_0639_),
    .A2(_0811_),
    .ZN(_0868_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4194_ (.A1(_0644_),
    .A2(_0804_),
    .ZN(_0869_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4195_ (.A1(_0638_),
    .A2(_0805_),
    .B1(_0869_),
    .B2(_0810_),
    .ZN(_0870_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4196_ (.I(\mod.Arithmetic.CN.I_in[26] ),
    .Z(_0871_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _4197_ (.A1(\mod.Arithmetic.CN.I_in[24] ),
    .A2(_0871_),
    .A3(_0808_),
    .Z(_0872_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _4198_ (.A1(_0807_),
    .A2(\mod.Arithmetic.CN.I_in[26] ),
    .Z(_0873_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4199_ (.A1(\mod.Arithmetic.CN.I_in[24] ),
    .A2(_0809_),
    .B(_0873_),
    .ZN(_0874_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4200_ (.A1(_0844_),
    .A2(\mod.Arithmetic.CN.I_in[18] ),
    .ZN(_0875_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _4201_ (.A1(_0803_),
    .A2(_0875_),
    .ZN(_0876_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4202_ (.A1(_0872_),
    .A2(_0874_),
    .B(_0876_),
    .ZN(_0877_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4203_ (.I(_0877_),
    .Z(_0878_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _4204_ (.A1(_0876_),
    .A2(_0872_),
    .A3(_0874_),
    .Z(_0879_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4205_ (.A1(_0878_),
    .A2(_0879_),
    .ZN(_0880_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _4206_ (.A1(_0868_),
    .A2(_0870_),
    .A3(_0880_),
    .Z(_0881_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4207_ (.A1(_0813_),
    .A2(_0715_),
    .ZN(_0882_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4208_ (.A1(\mod.Arithmetic.CN.I_in[8] ),
    .A2(_0814_),
    .B(_0882_),
    .ZN(_0883_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _4209_ (.A1(\mod.Arithmetic.CN.I_in[8] ),
    .A2(_0707_),
    .A3(_0814_),
    .B(_0883_),
    .ZN(_0884_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _4210_ (.A1(_0881_),
    .A2(_0884_),
    .ZN(_0885_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4211_ (.A1(_0867_),
    .A2(_0885_),
    .Z(_0886_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4212_ (.A1(_0825_),
    .A2(_0849_),
    .ZN(_0887_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4213_ (.A1(_0825_),
    .A2(_0849_),
    .ZN(_0888_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4214_ (.A1(_0836_),
    .A2(_0887_),
    .B(_0888_),
    .ZN(_0889_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4215_ (.A1(_0830_),
    .A2(_0834_),
    .ZN(_0890_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4216_ (.I(_0653_),
    .Z(_0891_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _4217_ (.A1(_0891_),
    .A2(\mod.Arithmetic.CN.I_in[34] ),
    .ZN(_0892_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4218_ (.I(\mod.Arithmetic.CN.I_in[34] ),
    .Z(_0893_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4219_ (.A1(_0820_),
    .A2(_0826_),
    .ZN(_0894_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _4220_ (.I0(_0892_),
    .I1(_0893_),
    .S(_0894_),
    .Z(_0895_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4221_ (.A1(_0643_),
    .A2(\mod.Arithmetic.CN.I_in[42] ),
    .ZN(_0896_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4222_ (.I(\mod.Arithmetic.CN.I_in[42] ),
    .Z(_0897_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4223_ (.A1(_0656_),
    .A2(_0831_),
    .ZN(_0898_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _4224_ (.I0(_0896_),
    .I1(_0897_),
    .S(_0898_),
    .Z(_0899_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4225_ (.A1(_0895_),
    .A2(_0899_),
    .Z(_0900_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _4226_ (.A1(_0890_),
    .A2(_0900_),
    .Z(_0901_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4227_ (.A1(_0890_),
    .A2(_0900_),
    .ZN(_0902_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4228_ (.A1(_0901_),
    .A2(_0902_),
    .ZN(_0903_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4229_ (.I(_0839_),
    .ZN(_0904_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _4230_ (.A1(_0837_),
    .A2(_0848_),
    .Z(_0905_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _4231_ (.A1(_0837_),
    .A2(_0848_),
    .Z(_0906_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4232_ (.A1(_0904_),
    .A2(_0905_),
    .B(_0906_),
    .ZN(_0907_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4233_ (.A1(_0662_),
    .A2(_0847_),
    .Z(_0908_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _4234_ (.A1(_0619_),
    .A2(_0661_),
    .A3(\mod.Arithmetic.CN.I_in[64] ),
    .A4(_0847_),
    .ZN(_0909_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4235_ (.A1(_0841_),
    .A2(_0908_),
    .B(_0909_),
    .ZN(_0910_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4236_ (.A1(_0664_),
    .A2(_0846_),
    .ZN(_0911_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _4237_ (.A1(_0665_),
    .A2(_0846_),
    .Z(_0912_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _4238_ (.A1(_0842_),
    .A2(_0911_),
    .A3(_0912_),
    .Z(_0913_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _4239_ (.A1(_0615_),
    .A2(\mod.Arithmetic.CN.I_in[66] ),
    .ZN(_0914_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4240_ (.I(_0807_),
    .Z(_0915_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _4241_ (.A1(_0915_),
    .A2(\mod.Arithmetic.ACTI.x[1] ),
    .A3(_0663_),
    .ZN(_0916_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4242_ (.A1(_0615_),
    .A2(\mod.Arithmetic.ACTI.x[2] ),
    .ZN(_0917_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4243_ (.A1(_0842_),
    .A2(_0917_),
    .Z(_0918_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4244_ (.A1(_0916_),
    .A2(_0918_),
    .Z(_0919_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _4245_ (.A1(_0911_),
    .A2(_0914_),
    .A3(_0919_),
    .ZN(_0920_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4246_ (.A1(_0913_),
    .A2(_0920_),
    .Z(_0921_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4247_ (.I(\mod.Arithmetic.CN.I_in[58] ),
    .Z(_0922_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4248_ (.I(_0922_),
    .Z(_0923_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _4249_ (.A1(_0619_),
    .A2(\mod.Arithmetic.CN.I_in[57] ),
    .A3(_0660_),
    .ZN(_0924_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _4250_ (.A1(_0637_),
    .A2(_0922_),
    .A3(_0924_),
    .ZN(_0925_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _4251_ (.A1(_0923_),
    .A2(_0924_),
    .B(_0925_),
    .ZN(_0926_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _4252_ (.A1(_0910_),
    .A2(_0921_),
    .A3(_0926_),
    .Z(_0927_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4253_ (.I(\mod.Arithmetic.CN.I_in[50] ),
    .Z(_0928_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4254_ (.I(_0928_),
    .Z(_0929_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4255_ (.I(\mod.Arithmetic.CN.I_in[49] ),
    .Z(_0930_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _4256_ (.A1(_0621_),
    .A2(_0930_),
    .A3(_0658_),
    .ZN(_0931_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _4257_ (.A1(_0824_),
    .A2(_0929_),
    .A3(_0931_),
    .ZN(_0932_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _4258_ (.A1(_0929_),
    .A2(_0931_),
    .B(_0932_),
    .ZN(_0933_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _4259_ (.A1(_0907_),
    .A2(_0927_),
    .A3(_0933_),
    .Z(_0934_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _4260_ (.A1(_0889_),
    .A2(_0903_),
    .A3(_0934_),
    .ZN(_0935_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _4261_ (.A1(_0866_),
    .A2(_0886_),
    .A3(_0935_),
    .ZN(_0936_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4262_ (.A1(_0865_),
    .A2(_0936_),
    .Z(_0937_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4263_ (.A1(_0862_),
    .A2(_0937_),
    .Z(_0938_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _4264_ (.A1(_0861_),
    .A2(_0938_),
    .ZN(_0939_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _4265_ (.I0(_0768_),
    .I1(_0773_),
    .S(_0794_),
    .Z(_0940_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _4266_ (.A1(_0768_),
    .A2(_0855_),
    .B1(_0857_),
    .B2(_0940_),
    .C(_0627_),
    .ZN(_0941_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4267_ (.A1(_0629_),
    .A2(_0939_),
    .B(_0941_),
    .ZN(\mod.P3.Res[2] ));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4268_ (.A1(_0861_),
    .A2(_0938_),
    .ZN(_0942_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4269_ (.I(_0862_),
    .ZN(_0943_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _4270_ (.A1(_0865_),
    .A2(_0936_),
    .Z(_0944_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4271_ (.A1(_0943_),
    .A2(_0937_),
    .B(_0944_),
    .ZN(_0945_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4272_ (.A1(_0867_),
    .A2(_0885_),
    .ZN(_0946_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _4273_ (.A1(_0866_),
    .A2(_0886_),
    .Z(_0947_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4274_ (.A1(_0946_),
    .A2(_0947_),
    .ZN(_0948_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4275_ (.A1(_0866_),
    .A2(_0886_),
    .ZN(_0949_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4276_ (.A1(_0903_),
    .A2(_0934_),
    .Z(_0950_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _4277_ (.A1(_0947_),
    .A2(_0949_),
    .A3(_0935_),
    .B1(_0950_),
    .B2(_0889_),
    .ZN(_0951_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4278_ (.A1(_0881_),
    .A2(_0884_),
    .ZN(_0952_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4279_ (.A1(_0687_),
    .A2(_0804_),
    .ZN(_0953_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _4280_ (.A1(_0871_),
    .A2(_0646_),
    .A3(_0809_),
    .ZN(_0954_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4281_ (.A1(_0877_),
    .A2(_0954_),
    .ZN(_0955_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4282_ (.A1(_0806_),
    .A2(\mod.Arithmetic.CN.I_in[19] ),
    .ZN(_0956_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _4283_ (.A1(_0875_),
    .A2(_0956_),
    .ZN(_0957_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4284_ (.I(\mod.Arithmetic.CN.I_in[27] ),
    .Z(_0958_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4285_ (.I(_0958_),
    .Z(_0959_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _4286_ (.A1(_0959_),
    .A2(_0808_),
    .A3(_0873_),
    .Z(_0960_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _4287_ (.A1(_0915_),
    .A2(_0959_),
    .B1(_0808_),
    .B2(_0873_),
    .ZN(_0961_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _4288_ (.A1(_0957_),
    .A2(_0960_),
    .A3(_0961_),
    .Z(_0962_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4289_ (.A1(_0960_),
    .A2(_0961_),
    .B(_0957_),
    .ZN(_0963_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _4290_ (.A1(_0962_),
    .A2(_0963_),
    .Z(_0964_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _4291_ (.A1(_0953_),
    .A2(_0955_),
    .A3(_0964_),
    .Z(_0965_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _4292_ (.A1(_0870_),
    .A2(_0878_),
    .A3(_0879_),
    .Z(_0966_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4293_ (.A1(_0878_),
    .A2(_0879_),
    .B(_0870_),
    .ZN(_0967_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _4294_ (.A1(_0868_),
    .A2(_0966_),
    .A3(_0967_),
    .ZN(_0968_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4295_ (.A1(_0966_),
    .A2(_0968_),
    .ZN(_0969_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4296_ (.A1(_0965_),
    .A2(_0969_),
    .Z(_0970_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4297_ (.A1(_0618_),
    .A2(\mod.Arithmetic.CN.I_in[11] ),
    .ZN(_0971_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4298_ (.I(_0971_),
    .Z(_0972_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _4299_ (.A1(_0716_),
    .A2(_0816_),
    .B1(_0882_),
    .B2(_0709_),
    .ZN(_0973_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4300_ (.A1(_0972_),
    .A2(_0973_),
    .Z(_0974_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _4301_ (.A1(_0901_),
    .A2(_0970_),
    .A3(_0974_),
    .Z(_0975_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _4302_ (.A1(_0952_),
    .A2(_0975_),
    .ZN(_0976_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _4303_ (.A1(_0927_),
    .A2(_0933_),
    .ZN(_0977_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _4304_ (.A1(_0901_),
    .A2(_0902_),
    .A3(_0934_),
    .B1(_0977_),
    .B2(_0907_),
    .ZN(_0978_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _4305_ (.A1(_0895_),
    .A2(_0899_),
    .Z(_0979_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _4306_ (.A1(_0891_),
    .A2(\mod.Arithmetic.CN.I_in[35] ),
    .ZN(_0980_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _4307_ (.A1(_0893_),
    .A2(_0829_),
    .B1(_0892_),
    .B2(\mod.Arithmetic.CN.I_in[33] ),
    .ZN(_0981_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _4308_ (.A1(_0980_),
    .A2(_0981_),
    .ZN(_0982_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4309_ (.A1(_0650_),
    .A2(\mod.Arithmetic.CN.I_in[43] ),
    .ZN(_0983_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4310_ (.I(_0983_),
    .Z(_0984_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _4311_ (.A1(_0897_),
    .A2(_0833_),
    .B1(_0896_),
    .B2(\mod.Arithmetic.CN.I_in[41] ),
    .ZN(_0985_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4312_ (.A1(_0984_),
    .A2(_0985_),
    .Z(_0986_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4313_ (.A1(_0982_),
    .A2(_0986_),
    .Z(_0987_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _4314_ (.A1(_0979_),
    .A2(_0987_),
    .ZN(_0988_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _4315_ (.A1(_0979_),
    .A2(_0987_),
    .Z(_0989_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _4316_ (.A1(_0988_),
    .A2(_0989_),
    .Z(_0990_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4317_ (.A1(_0921_),
    .A2(_0926_),
    .Z(_0991_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4318_ (.A1(_0910_),
    .A2(_0991_),
    .B1(_0927_),
    .B2(_0933_),
    .ZN(_0992_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _4319_ (.A1(_0929_),
    .A2(_0658_),
    .A3(_0838_),
    .ZN(_0993_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _4320_ (.A1(_0922_),
    .A2(_0660_),
    .A3(_0840_),
    .ZN(_0994_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _4321_ (.A1(_0654_),
    .A2(_0928_),
    .A3(\mod.Arithmetic.CN.I_in[51] ),
    .ZN(_0995_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _4322_ (.A1(_0891_),
    .A2(\mod.Arithmetic.CN.I_in[50] ),
    .A3(_0838_),
    .Z(_0996_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _4323_ (.A1(_0653_),
    .A2(\mod.Arithmetic.CN.I_in[51] ),
    .Z(_0997_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _4324_ (.A1(_0930_),
    .A2(_0995_),
    .B1(_0996_),
    .B2(_0997_),
    .ZN(_0998_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _4325_ (.A1(_0994_),
    .A2(_0998_),
    .ZN(_0999_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _4326_ (.A1(_0993_),
    .A2(_0999_),
    .Z(_1000_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4327_ (.A1(_0993_),
    .A2(_0999_),
    .ZN(_1001_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4328_ (.A1(_1000_),
    .A2(_1001_),
    .ZN(_1002_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4329_ (.A1(_0913_),
    .A2(_0920_),
    .ZN(_1003_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _4330_ (.A1(_0921_),
    .A2(_0926_),
    .B(_1003_),
    .ZN(_1004_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4331_ (.A1(_0911_),
    .A2(_0919_),
    .Z(_1005_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _4332_ (.A1(_0665_),
    .A2(_0846_),
    .A3(_0919_),
    .Z(_1006_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _4333_ (.A1(_0914_),
    .A2(_1005_),
    .B(_1006_),
    .ZN(_1007_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _4334_ (.A1(_0640_),
    .A2(\mod.Arithmetic.CN.I_in[67] ),
    .Z(_1008_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _4335_ (.A1(\mod.Arithmetic.CN.I_in[64] ),
    .A2(_0918_),
    .B(\mod.Arithmetic.ACTI.x[1] ),
    .C(_0643_),
    .ZN(_1009_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _4336_ (.A1(_0642_),
    .A2(\mod.Arithmetic.ACTI.x[2] ),
    .A3(_0842_),
    .ZN(_1010_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4337_ (.A1(_0641_),
    .A2(\mod.Arithmetic.ACTI.x[3] ),
    .ZN(_1011_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4338_ (.A1(_0914_),
    .A2(_1011_),
    .Z(_1012_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4339_ (.A1(_1010_),
    .A2(_1012_),
    .Z(_1013_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4340_ (.A1(_1009_),
    .A2(_1013_),
    .Z(_1014_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4341_ (.A1(_1008_),
    .A2(_1014_),
    .Z(_1015_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4342_ (.A1(_1007_),
    .A2(_1015_),
    .Z(_1016_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4343_ (.I(\mod.Arithmetic.CN.I_in[59] ),
    .Z(_1017_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4344_ (.I(_1017_),
    .Z(_1018_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4345_ (.A1(_0617_),
    .A2(_1017_),
    .ZN(_1019_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _4346_ (.A1(_0813_),
    .A2(_0923_),
    .A3(_0840_),
    .ZN(_1020_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _4347_ (.I0(_1018_),
    .I1(_1019_),
    .S(_1020_),
    .Z(_1021_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _4348_ (.A1(_1004_),
    .A2(_1016_),
    .A3(_1021_),
    .Z(_1022_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _4349_ (.A1(_0992_),
    .A2(_1002_),
    .A3(_1022_),
    .Z(_1023_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _4350_ (.A1(_0978_),
    .A2(_0990_),
    .A3(_1023_),
    .ZN(_1024_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _4351_ (.A1(_0951_),
    .A2(_0976_),
    .A3(_1024_),
    .ZN(_1025_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _4352_ (.A1(_0948_),
    .A2(_1025_),
    .ZN(_1026_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _4353_ (.A1(_0945_),
    .A2(_1026_),
    .ZN(_1027_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4354_ (.A1(_0942_),
    .A2(_1027_),
    .Z(_1028_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _4355_ (.I0(_0775_),
    .I1(_0774_),
    .S(_0794_),
    .Z(_1029_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _4356_ (.A1(_0775_),
    .A2(_0855_),
    .B1(_0856_),
    .B2(_1029_),
    .C(_0627_),
    .ZN(_1030_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4357_ (.A1(_0629_),
    .A2(_1028_),
    .B(_1030_),
    .ZN(\mod.P3.Res[3] ));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4358_ (.I(_0627_),
    .Z(_1031_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4359_ (.A1(_0781_),
    .A2(_0799_),
    .ZN(_1032_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4360_ (.A1(_0780_),
    .A2(_0795_),
    .ZN(_1033_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4361_ (.A1(_0781_),
    .A2(_0854_),
    .B1(_0856_),
    .B2(_1033_),
    .ZN(_1034_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4362_ (.A1(_0945_),
    .A2(_1026_),
    .ZN(_1035_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _4363_ (.A1(_0861_),
    .A2(_0938_),
    .A3(_1027_),
    .ZN(_1036_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4364_ (.A1(_0976_),
    .A2(_1024_),
    .Z(_1037_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4365_ (.A1(_0948_),
    .A2(_1025_),
    .ZN(_1038_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4366_ (.A1(_0951_),
    .A2(_1037_),
    .B(_1038_),
    .ZN(_1039_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4367_ (.A1(_0970_),
    .A2(_0974_),
    .Z(_1040_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _4368_ (.A1(_0901_),
    .A2(_1040_),
    .Z(_1041_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4369_ (.A1(_0952_),
    .A2(_0975_),
    .B(_1041_),
    .ZN(_1042_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4370_ (.A1(_0990_),
    .A2(_1023_),
    .Z(_1043_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _4371_ (.A1(_0978_),
    .A2(_1043_),
    .Z(_1044_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4372_ (.A1(_0976_),
    .A2(_1024_),
    .ZN(_1045_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4373_ (.A1(_1044_),
    .A2(_1045_),
    .ZN(_1046_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4374_ (.A1(_0970_),
    .A2(_0974_),
    .ZN(_1047_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4375_ (.A1(_0968_),
    .A2(_0965_),
    .ZN(_1048_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4376_ (.A1(_0966_),
    .A2(_0965_),
    .ZN(_1049_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _4377_ (.A1(_0962_),
    .A2(_0963_),
    .B(_0877_),
    .C(_0954_),
    .ZN(_1050_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4378_ (.A1(_0878_),
    .A2(_0954_),
    .B(_0962_),
    .C(_0963_),
    .ZN(_1051_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _4379_ (.A1(_0687_),
    .A2(_0804_),
    .A3(_1050_),
    .B(_1051_),
    .ZN(_1052_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _4380_ (.A1(_0617_),
    .A2(_0680_),
    .A3(_0682_),
    .ZN(_1053_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _4381_ (.A1(_0957_),
    .A2(_0960_),
    .A3(_0961_),
    .ZN(_1054_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _4382_ (.A1(_0844_),
    .A2(\mod.Arithmetic.CN.I_in[26] ),
    .ZN(_1055_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _4383_ (.A1(_0634_),
    .A2(_0959_),
    .B(_0809_),
    .C(_1055_),
    .ZN(_1056_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4384_ (.A1(_1054_),
    .A2(_1056_),
    .ZN(_1057_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _4385_ (.A1(_0616_),
    .A2(_0691_),
    .A3(\mod.Arithmetic.CN.I_in[19] ),
    .ZN(_1058_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4386_ (.A1(_0806_),
    .A2(\mod.Arithmetic.CN.I_in[20] ),
    .ZN(_1059_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4387_ (.A1(_0956_),
    .A2(_1059_),
    .ZN(_1060_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4388_ (.I(_0632_),
    .ZN(_1061_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4389_ (.I(\mod.Arithmetic.CN.I_in[28] ),
    .Z(_1062_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4390_ (.I(_1062_),
    .ZN(_1063_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4391_ (.A1(_0843_),
    .A2(\mod.Arithmetic.CN.I_in[27] ),
    .ZN(_1064_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _4392_ (.A1(_1061_),
    .A2(_1063_),
    .B1(_1064_),
    .B2(_0871_),
    .ZN(_1065_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _4393_ (.A1(_0642_),
    .A2(_0959_),
    .A3(_1062_),
    .A4(_1055_),
    .ZN(_1066_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _4394_ (.A1(_1058_),
    .A2(_1060_),
    .A3(_1065_),
    .A4(_1066_),
    .ZN(_1067_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _4395_ (.A1(_0956_),
    .A2(_1059_),
    .ZN(_1068_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _4396_ (.A1(_0615_),
    .A2(_0958_),
    .A3(_1063_),
    .A4(_1055_),
    .ZN(_1069_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _4397_ (.A1(_0843_),
    .A2(\mod.Arithmetic.CN.I_in[28] ),
    .Z(_1070_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4398_ (.A1(_0871_),
    .A2(_1064_),
    .B(_1070_),
    .ZN(_1071_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _4399_ (.A1(_1068_),
    .A2(_1069_),
    .A3(_1071_),
    .ZN(_1072_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4400_ (.A1(_1067_),
    .A2(_1072_),
    .ZN(_1073_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _4401_ (.A1(_1053_),
    .A2(_1057_),
    .A3(_1073_),
    .ZN(_1074_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4402_ (.A1(_1052_),
    .A2(_1074_),
    .Z(_1075_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _4403_ (.A1(_0893_),
    .A2(_0829_),
    .A3(_0980_),
    .ZN(_1076_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _4404_ (.A1(_1049_),
    .A2(_1075_),
    .A3(_1076_),
    .Z(_1077_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4405_ (.A1(_0620_),
    .A2(_0724_),
    .ZN(_1078_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _4406_ (.A1(_0813_),
    .A2(_0722_),
    .A3(_0715_),
    .A4(\mod.Arithmetic.CN.I_in[9] ),
    .ZN(_1079_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4407_ (.A1(_0715_),
    .A2(_0972_),
    .B(_1079_),
    .ZN(_1080_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _4408_ (.A1(_0716_),
    .A2(_0816_),
    .A3(_0972_),
    .B(_1080_),
    .ZN(_1081_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4409_ (.A1(_1078_),
    .A2(_1081_),
    .Z(_1082_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _4410_ (.A1(_1048_),
    .A2(_1077_),
    .A3(_1082_),
    .Z(_1083_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4411_ (.A1(_0988_),
    .A2(_1083_),
    .Z(_1084_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _4412_ (.A1(_1002_),
    .A2(_1022_),
    .Z(_1085_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4413_ (.A1(_1002_),
    .A2(_1022_),
    .ZN(_1086_));
 gf180mcu_fd_sc_mcu7t5v0__oai33_1 _4414_ (.A1(_0992_),
    .A2(_1085_),
    .A3(_1086_),
    .B1(_1023_),
    .B2(_0988_),
    .B3(_0989_),
    .ZN(_1087_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4415_ (.I(_0986_),
    .ZN(_1088_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4416_ (.A1(_0982_),
    .A2(_1088_),
    .ZN(_1089_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4417_ (.I(\mod.Arithmetic.CN.I_in[36] ),
    .Z(_1090_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4418_ (.A1(_0655_),
    .A2(_1090_),
    .ZN(_1091_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4419_ (.A1(_0893_),
    .A2(_0980_),
    .ZN(_1092_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_4 _4420_ (.A1(_0828_),
    .A2(\mod.Arithmetic.CN.I_in[35] ),
    .B(_0826_),
    .C(_0892_),
    .ZN(_1093_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4421_ (.A1(_1092_),
    .A2(_1093_),
    .ZN(_1094_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4422_ (.A1(_1091_),
    .A2(_1094_),
    .Z(_1095_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4423_ (.A1(_0654_),
    .A2(\mod.Arithmetic.CN.I_in[44] ),
    .ZN(_1096_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _4424_ (.A1(_0897_),
    .A2(_0984_),
    .Z(_1097_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _4425_ (.A1(_0619_),
    .A2(\mod.Arithmetic.CN.I_in[41] ),
    .A3(_0897_),
    .A4(_0984_),
    .ZN(_1098_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4426_ (.A1(_0833_),
    .A2(_1097_),
    .ZN(_1099_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4427_ (.A1(_1097_),
    .A2(_1098_),
    .B(_1099_),
    .ZN(_1100_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4428_ (.A1(_1096_),
    .A2(_1100_),
    .Z(_1101_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4429_ (.A1(_1095_),
    .A2(_1101_),
    .Z(_1102_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4430_ (.A1(_1089_),
    .A2(_1102_),
    .Z(_1103_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _4431_ (.A1(_0824_),
    .A2(_1018_),
    .A3(_1020_),
    .ZN(_1104_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4432_ (.A1(_1018_),
    .A2(_1020_),
    .B(_1104_),
    .ZN(_1105_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _4433_ (.A1(_1004_),
    .A2(_1016_),
    .A3(_1105_),
    .Z(_1106_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4434_ (.A1(_1016_),
    .A2(_1021_),
    .Z(_1107_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_2 _4435_ (.A1(_1000_),
    .A2(_1001_),
    .A3(_1106_),
    .B1(_1107_),
    .B2(_1004_),
    .ZN(_1108_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _4436_ (.A1(_0930_),
    .A2(_0995_),
    .B1(_0996_),
    .B2(_0997_),
    .C(_0994_),
    .ZN(_1109_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4437_ (.A1(_0993_),
    .A2(_0999_),
    .ZN(_1110_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4438_ (.A1(_1109_),
    .A2(_1110_),
    .ZN(_1111_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _4439_ (.A1(_0650_),
    .A2(\mod.Arithmetic.CN.I_in[57] ),
    .A3(_0922_),
    .A4(_1019_),
    .Z(_1112_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4440_ (.A1(\mod.Arithmetic.CN.I_in[52] ),
    .A2(_0997_),
    .ZN(_1113_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4441_ (.A1(_0616_),
    .A2(\mod.Arithmetic.CN.I_in[51] ),
    .ZN(_1114_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4442_ (.A1(\mod.Arithmetic.CN.I_in[50] ),
    .A2(_1114_),
    .ZN(_1115_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _4443_ (.A1(_0915_),
    .A2(\mod.Arithmetic.CN.I_in[52] ),
    .Z(_1116_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _4444_ (.A1(_0928_),
    .A2(_1113_),
    .B1(_1115_),
    .B2(_1116_),
    .ZN(_1117_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4445_ (.A1(_1112_),
    .A2(_1117_),
    .Z(_1118_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _4446_ (.A1(_0828_),
    .A2(_0930_),
    .A3(_0928_),
    .A4(_1114_),
    .ZN(_1119_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4447_ (.A1(_1118_),
    .A2(_1119_),
    .Z(_1120_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4448_ (.A1(_1111_),
    .A2(_1120_),
    .Z(_1121_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _4449_ (.A1(_1007_),
    .A2(_1015_),
    .B1(_1016_),
    .B2(_1105_),
    .ZN(_1122_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4450_ (.A1(_1009_),
    .A2(_1013_),
    .ZN(_1123_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4451_ (.A1(_1008_),
    .A2(_1014_),
    .B(_1123_),
    .ZN(_1124_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4452_ (.A1(_0614_),
    .A2(\mod.Arithmetic.CN.I_in[68] ),
    .ZN(_1125_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _4453_ (.A1(\mod.Arithmetic.CN.I_in[65] ),
    .A2(_1012_),
    .B(_0645_),
    .C(\mod.Arithmetic.ACTI.x[2] ),
    .ZN(_1126_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _4454_ (.A1(_0915_),
    .A2(\mod.Arithmetic.ACTI.x[3] ),
    .A3(_0914_),
    .ZN(_1127_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4455_ (.A1(_0640_),
    .A2(\mod.Arithmetic.ACTI.x[4] ),
    .ZN(_1128_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _4456_ (.A1(_1008_),
    .A2(_1128_),
    .ZN(_1129_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4457_ (.A1(_1127_),
    .A2(_1129_),
    .Z(_1130_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4458_ (.A1(_1126_),
    .A2(_1130_),
    .Z(_1131_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4459_ (.A1(_1125_),
    .A2(_1131_),
    .Z(_1132_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _4460_ (.A1(_1124_),
    .A2(_1132_),
    .ZN(_1133_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4461_ (.I(\mod.Arithmetic.CN.I_in[60] ),
    .Z(_1134_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _4462_ (.A1(_0635_),
    .A2(_1017_),
    .A3(_1134_),
    .ZN(_1135_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4463_ (.A1(_0642_),
    .A2(\mod.Arithmetic.CN.I_in[60] ),
    .ZN(_1136_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4464_ (.A1(_0923_),
    .A2(_1019_),
    .B(_1136_),
    .ZN(_1137_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4465_ (.A1(_0923_),
    .A2(_1135_),
    .B(_1137_),
    .ZN(_1138_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _4466_ (.A1(_1133_),
    .A2(_1138_),
    .ZN(_1139_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _4467_ (.A1(_1121_),
    .A2(_1122_),
    .A3(_1139_),
    .Z(_1140_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _4468_ (.A1(_1103_),
    .A2(_1108_),
    .A3(_1140_),
    .Z(_1141_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4469_ (.A1(_1087_),
    .A2(_1141_),
    .Z(_1142_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _4470_ (.A1(_1047_),
    .A2(_1084_),
    .A3(_1142_),
    .Z(_1143_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _4471_ (.A1(_1042_),
    .A2(_1046_),
    .A3(_1143_),
    .ZN(_1144_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4472_ (.A1(_1039_),
    .A2(_1144_),
    .Z(_1145_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _4473_ (.A1(_1035_),
    .A2(_1036_),
    .A3(_1145_),
    .Z(_1146_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4474_ (.A1(_1035_),
    .A2(_1036_),
    .B(_1145_),
    .ZN(_1147_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _4475_ (.A1(_1031_),
    .A2(_1146_),
    .A3(_1147_),
    .ZN(_1148_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _4476_ (.A1(_1031_),
    .A2(_1032_),
    .A3(_1034_),
    .B(_1148_),
    .ZN(\mod.P3.Res[4] ));
 gf180mcu_fd_sc_mcu7t5v0__nor4_2 _4477_ (.A1(_0725_),
    .A2(_0716_),
    .A3(_0816_),
    .A4(_0972_),
    .ZN(_1149_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _4478_ (.A1(_1044_),
    .A2(_1045_),
    .A3(_1143_),
    .ZN(_1150_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4479_ (.A1(_1044_),
    .A2(_1045_),
    .B(_1143_),
    .ZN(_1151_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4480_ (.A1(_1042_),
    .A2(_1150_),
    .B(_1151_),
    .ZN(_1152_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _4481_ (.A1(_1047_),
    .A2(_1084_),
    .Z(_1153_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4482_ (.A1(_0988_),
    .A2(_1083_),
    .B(_1153_),
    .ZN(_1154_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4483_ (.A1(_1047_),
    .A2(_1084_),
    .ZN(_1155_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4484_ (.A1(_1087_),
    .A2(_1141_),
    .ZN(_1156_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4485_ (.A1(_1087_),
    .A2(_1141_),
    .ZN(_1157_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _4486_ (.A1(_1153_),
    .A2(_1155_),
    .A3(_1156_),
    .B(_1157_),
    .ZN(_1158_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4487_ (.A1(_1089_),
    .A2(_1102_),
    .ZN(_1159_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _4488_ (.A1(_1048_),
    .A2(_1077_),
    .Z(_1160_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _4489_ (.A1(_1048_),
    .A2(_1077_),
    .Z(_1161_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4490_ (.A1(_1160_),
    .A2(_1082_),
    .B(_1161_),
    .ZN(_1162_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _4491_ (.A1(_1075_),
    .A2(_1076_),
    .Z(_1163_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _4492_ (.A1(_1075_),
    .A2(_1076_),
    .Z(_1164_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4493_ (.A1(_1049_),
    .A2(_1163_),
    .B(_1164_),
    .ZN(_1165_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4494_ (.A1(_1052_),
    .A2(_1074_),
    .ZN(_1166_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _4495_ (.A1(_1067_),
    .A2(_1072_),
    .B(_1054_),
    .C(_1056_),
    .ZN(_1167_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4496_ (.A1(_1054_),
    .A2(_1056_),
    .B(_1067_),
    .C(_1072_),
    .ZN(_1168_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4497_ (.A1(_1053_),
    .A2(_1167_),
    .B(_1168_),
    .ZN(_1169_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4498_ (.A1(_1069_),
    .A2(_1071_),
    .B(_1068_),
    .ZN(_1170_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _4499_ (.A1(_1055_),
    .A2(_1064_),
    .A3(_1070_),
    .ZN(_1171_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4500_ (.A1(_1170_),
    .A2(_1171_),
    .ZN(_1172_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4501_ (.A1(_0678_),
    .A2(\mod.Arithmetic.CN.I_in[20] ),
    .B(_0843_),
    .ZN(_1173_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _4502_ (.A1(_0613_),
    .A2(\mod.Arithmetic.CN.I_in[21] ),
    .A3(\mod.Arithmetic.CN.I_in[20] ),
    .Z(_1174_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _4503_ (.A1(_1173_),
    .A2(_1174_),
    .Z(_1175_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _4504_ (.A1(_0806_),
    .A2(_1062_),
    .A3(\mod.Arithmetic.CN.I_in[29] ),
    .ZN(_1176_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4505_ (.A1(_0958_),
    .A2(_1176_),
    .ZN(_1177_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4506_ (.I(\mod.Arithmetic.CN.I_in[29] ),
    .Z(_1178_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4507_ (.A1(_0632_),
    .A2(_1178_),
    .B1(_1064_),
    .B2(_1070_),
    .ZN(_1179_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _4508_ (.A1(_1175_),
    .A2(_1177_),
    .A3(_1179_),
    .Z(_1180_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4509_ (.A1(_1177_),
    .A2(_1179_),
    .B(_1175_),
    .ZN(_1181_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4510_ (.A1(_1180_),
    .A2(_1181_),
    .ZN(_1182_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _4511_ (.A1(_1058_),
    .A2(_1172_),
    .A3(_1182_),
    .ZN(_1183_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4512_ (.A1(_1169_),
    .A2(_1183_),
    .Z(_1184_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4513_ (.I(_1090_),
    .Z(_1185_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4514_ (.A1(_1185_),
    .A2(_1093_),
    .ZN(_1186_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _4515_ (.A1(_1166_),
    .A2(_1184_),
    .A3(_1186_),
    .ZN(_1187_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4516_ (.A1(_0824_),
    .A2(_0731_),
    .ZN(_1188_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4517_ (.I(\mod.Arithmetic.CN.I_in[12] ),
    .ZN(_1189_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4518_ (.I(_1189_),
    .Z(_1190_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _4519_ (.A1(_0724_),
    .A2(_0707_),
    .A3(_0971_),
    .ZN(_1191_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4520_ (.A1(\mod.Arithmetic.CN.I_in[11] ),
    .A2(_1078_),
    .ZN(_1192_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _4521_ (.A1(_1190_),
    .A2(_1079_),
    .B1(_1191_),
    .B2(_1192_),
    .ZN(_1193_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _4522_ (.A1(_1188_),
    .A2(_1193_),
    .ZN(_1194_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4523_ (.I(_1194_),
    .ZN(_1195_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _4524_ (.A1(_1165_),
    .A2(_1187_),
    .A3(_1195_),
    .Z(_1196_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _4525_ (.A1(_1159_),
    .A2(_1162_),
    .A3(_1196_),
    .Z(_1197_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4526_ (.I(_1103_),
    .ZN(_1198_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4527_ (.A1(_1108_),
    .A2(_1140_),
    .ZN(_1199_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4528_ (.A1(_1108_),
    .A2(_1140_),
    .ZN(_1200_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4529_ (.A1(_1198_),
    .A2(_1199_),
    .B(_1200_),
    .ZN(_1201_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4530_ (.I(\mod.Arithmetic.CN.I_in[44] ),
    .ZN(_1202_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4531_ (.I(_1202_),
    .Z(_1203_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4532_ (.I(_1101_),
    .ZN(_1204_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4533_ (.A1(_1203_),
    .A2(_1099_),
    .B1(_1204_),
    .B2(_1095_),
    .ZN(_1205_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _4534_ (.A1(_1203_),
    .A2(_1098_),
    .Z(_1206_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4535_ (.I(_1206_),
    .ZN(_1207_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4536_ (.A1(_0651_),
    .A2(\mod.Arithmetic.CN.I_in[45] ),
    .ZN(_1208_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _4537_ (.A1(_0654_),
    .A2(\mod.Arithmetic.CN.I_in[44] ),
    .B(_0896_),
    .C(_0983_),
    .ZN(_1209_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4538_ (.A1(\mod.Arithmetic.CN.I_in[43] ),
    .A2(_1096_),
    .ZN(_1210_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4539_ (.A1(_1209_),
    .A2(_1210_),
    .ZN(_1211_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _4540_ (.A1(_1208_),
    .A2(_1211_),
    .ZN(_1212_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4541_ (.A1(_0637_),
    .A2(\mod.Arithmetic.CN.I_in[37] ),
    .ZN(_1213_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _4542_ (.A1(_0636_),
    .A2(\mod.Arithmetic.CN.I_in[36] ),
    .B(_0892_),
    .C(_0980_),
    .ZN(_1214_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4543_ (.A1(\mod.Arithmetic.CN.I_in[35] ),
    .A2(_1091_),
    .ZN(_1215_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4544_ (.A1(_1214_),
    .A2(_1215_),
    .ZN(_1216_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4545_ (.A1(_1213_),
    .A2(_1216_),
    .Z(_1217_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _4546_ (.A1(_1207_),
    .A2(_1212_),
    .A3(_1217_),
    .Z(_1218_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _4547_ (.A1(_1205_),
    .A2(_1218_),
    .ZN(_1219_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4548_ (.A1(_1122_),
    .A2(_1139_),
    .ZN(_1220_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4549_ (.A1(_1122_),
    .A2(_1139_),
    .ZN(_1221_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4550_ (.A1(_1121_),
    .A2(_1220_),
    .B(_1221_),
    .ZN(_1222_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _4551_ (.A1(_0929_),
    .A2(_1113_),
    .B1(_1115_),
    .B2(_1116_),
    .C(_1112_),
    .ZN(_1223_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4552_ (.A1(_1118_),
    .A2(_1119_),
    .B(_1223_),
    .ZN(_1224_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4553_ (.I(\mod.Arithmetic.CN.I_in[52] ),
    .Z(_1225_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4554_ (.A1(_1225_),
    .A2(_0995_),
    .ZN(_1226_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _4555_ (.A1(_0653_),
    .A2(\mod.Arithmetic.CN.I_in[58] ),
    .A3(\mod.Arithmetic.CN.I_in[59] ),
    .A4(_1136_),
    .Z(_1227_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4556_ (.A1(_0645_),
    .A2(\mod.Arithmetic.CN.I_in[53] ),
    .B1(_1114_),
    .B2(_1116_),
    .ZN(_1228_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _4557_ (.A1(\mod.Arithmetic.CN.I_in[53] ),
    .A2(_1114_),
    .A3(_1116_),
    .Z(_1229_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4558_ (.A1(_1228_),
    .A2(_1229_),
    .ZN(_1230_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _4559_ (.A1(_1227_),
    .A2(_1230_),
    .ZN(_1231_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _4560_ (.A1(_1226_),
    .A2(_1231_),
    .ZN(_1232_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4561_ (.A1(_1224_),
    .A2(_1232_),
    .Z(_1233_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _4562_ (.A1(_1111_),
    .A2(_1120_),
    .A3(_1233_),
    .Z(_1234_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4563_ (.A1(_1111_),
    .A2(_1120_),
    .B(_1233_),
    .ZN(_1235_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _4564_ (.A1(_1234_),
    .A2(_1235_),
    .Z(_1236_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _4565_ (.A1(_1124_),
    .A2(_1132_),
    .B1(_1133_),
    .B2(_1138_),
    .ZN(_1237_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _4566_ (.A1(_0618_),
    .A2(\mod.Arithmetic.CN.I_in[68] ),
    .Z(_1238_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4567_ (.A1(_1126_),
    .A2(_1130_),
    .ZN(_1239_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4568_ (.A1(_1238_),
    .A2(_1131_),
    .B(_1239_),
    .ZN(_1240_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4569_ (.A1(_0614_),
    .A2(\mod.Arithmetic.CN.I_in[69] ),
    .ZN(_1241_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _4570_ (.A1(\mod.Arithmetic.CN.I_in[66] ),
    .A2(_1129_),
    .B(_0634_),
    .C(_0775_),
    .ZN(_1242_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4571_ (.A1(\mod.Arithmetic.CN.I_in[67] ),
    .A2(_1128_),
    .ZN(_1243_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4572_ (.A1(_0614_),
    .A2(\mod.Arithmetic.ACTI.x[5] ),
    .ZN(_1244_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4573_ (.A1(_1125_),
    .A2(_1244_),
    .Z(_1245_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _4574_ (.A1(_1243_),
    .A2(_1245_),
    .ZN(_1246_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4575_ (.A1(_1242_),
    .A2(_1246_),
    .Z(_1247_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4576_ (.A1(_1241_),
    .A2(_1247_),
    .Z(_1248_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _4577_ (.A1(_1240_),
    .A2(_1248_),
    .ZN(_1249_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4578_ (.I(\mod.Arithmetic.CN.I_in[61] ),
    .ZN(_1250_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4579_ (.I(_1061_),
    .Z(_1251_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _4580_ (.A1(_1251_),
    .A2(_1250_),
    .B1(_1136_),
    .B2(_1017_),
    .ZN(_1252_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _4581_ (.A1(_1018_),
    .A2(_1250_),
    .A3(_1136_),
    .B(_1252_),
    .ZN(_1253_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4582_ (.A1(_1249_),
    .A2(_1253_),
    .Z(_1254_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _4583_ (.A1(_1237_),
    .A2(_1254_),
    .ZN(_1255_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _4584_ (.A1(_1236_),
    .A2(_1255_),
    .ZN(_1256_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _4585_ (.A1(_1219_),
    .A2(_1222_),
    .A3(_1256_),
    .ZN(_1257_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _4586_ (.A1(_1197_),
    .A2(_1201_),
    .A3(_1257_),
    .ZN(_1258_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _4587_ (.A1(_1154_),
    .A2(_1158_),
    .A3(_1258_),
    .ZN(_1259_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _4588_ (.A1(_1149_),
    .A2(_1152_),
    .A3(_1259_),
    .Z(_1260_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4589_ (.A1(_1039_),
    .A2(_1144_),
    .B(_1147_),
    .ZN(_1261_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _4590_ (.A1(_1260_),
    .A2(_1261_),
    .ZN(_1262_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4591_ (.A1(_0785_),
    .A2(_0795_),
    .ZN(_1263_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4592_ (.A1(_0786_),
    .A2(_0799_),
    .B(_0857_),
    .C(_1263_),
    .ZN(_1264_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4593_ (.A1(_0786_),
    .A2(_0855_),
    .B(_0628_),
    .ZN(_1265_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4594_ (.A1(_1031_),
    .A2(_1262_),
    .B1(_1264_),
    .B2(_1265_),
    .ZN(\mod.P3.Res[5] ));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4595_ (.A1(_0799_),
    .A2(_0857_),
    .ZN(_1266_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _4596_ (.A1(\mod.P2.Rout_reg[0] ),
    .A2(_0672_),
    .Z(_1267_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _4597_ (.A1(\mod.Arithmetic.ACTI.x[6] ),
    .A2(_1267_),
    .A3(_0796_),
    .ZN(_1268_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4598_ (.A1(_1260_),
    .A2(_1261_),
    .ZN(_1269_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _4599_ (.A1(_1152_),
    .A2(_1259_),
    .Z(_1270_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _4600_ (.A1(_1152_),
    .A2(_1259_),
    .Z(_1271_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4601_ (.A1(_1149_),
    .A2(_1270_),
    .B(_1271_),
    .ZN(_1272_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _4602_ (.A1(_0625_),
    .A2(_0735_),
    .B(_1190_),
    .C(_1079_),
    .ZN(_1273_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4603_ (.A1(_1158_),
    .A2(_1258_),
    .ZN(_1274_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4604_ (.A1(_1158_),
    .A2(_1258_),
    .ZN(_1275_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4605_ (.A1(_1154_),
    .A2(_1274_),
    .B(_1275_),
    .ZN(_1276_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _4606_ (.A1(_1159_),
    .A2(_1196_),
    .ZN(_1277_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4607_ (.A1(_1162_),
    .A2(_1277_),
    .ZN(_1278_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4608_ (.A1(_1159_),
    .A2(_1196_),
    .B(_1278_),
    .ZN(_1279_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4609_ (.A1(_1201_),
    .A2(_1257_),
    .ZN(_1280_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4610_ (.A1(_1201_),
    .A2(_1257_),
    .ZN(_1281_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4611_ (.A1(_1197_),
    .A2(_1280_),
    .B(_1281_),
    .ZN(_1282_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4612_ (.A1(_1165_),
    .A2(_1187_),
    .ZN(_1283_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4613_ (.A1(_1165_),
    .A2(_1187_),
    .ZN(_1284_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4614_ (.A1(_1283_),
    .A2(_1195_),
    .B(_1284_),
    .ZN(_1285_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4615_ (.A1(_1205_),
    .A2(_1218_),
    .ZN(_1286_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4616_ (.I(\mod.Arithmetic.CN.I_in[13] ),
    .ZN(_1287_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4617_ (.I(\mod.Arithmetic.CN.I_in[14] ),
    .ZN(_1288_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4618_ (.A1(_1287_),
    .A2(_0724_),
    .B(_1288_),
    .ZN(_1289_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _4619_ (.A1(_0737_),
    .A2(\mod.Arithmetic.CN.I_in[13] ),
    .A3(_1190_),
    .ZN(_1290_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _4620_ (.A1(_0828_),
    .A2(_1289_),
    .A3(_1290_),
    .ZN(_1291_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4621_ (.A1(_0731_),
    .A2(_1191_),
    .ZN(_1292_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _4622_ (.A1(_1291_),
    .A2(_1292_),
    .Z(_1293_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _4623_ (.A1(\mod.Arithmetic.CN.I_in[13] ),
    .A2(_1189_),
    .A3(_0971_),
    .ZN(_1294_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _4624_ (.I0(_1291_),
    .I1(_0737_),
    .S(_1294_),
    .Z(_1295_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4625_ (.A1(_1292_),
    .A2(_1295_),
    .ZN(_1296_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4626_ (.A1(_1293_),
    .A2(_1296_),
    .ZN(_1297_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4627_ (.A1(_1185_),
    .A2(_1093_),
    .B(_1184_),
    .ZN(_1298_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _4628_ (.A1(_1185_),
    .A2(_1093_),
    .A3(_1184_),
    .ZN(_1299_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4629_ (.A1(_1166_),
    .A2(_1298_),
    .B(_1299_),
    .ZN(_1300_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4630_ (.A1(_1169_),
    .A2(_1183_),
    .ZN(_1301_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4631_ (.I(_1301_),
    .ZN(_1302_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4632_ (.A1(\mod.Arithmetic.CN.I_in[37] ),
    .A2(_1214_),
    .ZN(_1303_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _4633_ (.A1(_1180_),
    .A2(_1181_),
    .B(_1170_),
    .C(_1171_),
    .ZN(_1304_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4634_ (.A1(_1170_),
    .A2(_1171_),
    .B(_1180_),
    .C(_1181_),
    .ZN(_1305_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4635_ (.A1(_1058_),
    .A2(_1304_),
    .B(_1305_),
    .ZN(_1306_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4636_ (.I(_1178_),
    .ZN(_1307_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _4637_ (.A1(_0633_),
    .A2(_0958_),
    .A3(_1062_),
    .A4(_1307_),
    .ZN(_1308_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _4638_ (.A1(_1180_),
    .A2(_1308_),
    .Z(_1309_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _4639_ (.A1(_0844_),
    .A2(\mod.Arithmetic.CN.I_in[22] ),
    .A3(_0678_),
    .ZN(_1310_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4640_ (.A1(_0695_),
    .A2(_0679_),
    .B(_1061_),
    .ZN(_1311_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _4641_ (.A1(_1310_),
    .A2(_1311_),
    .Z(_1312_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _4642_ (.A1(_1063_),
    .A2(_1178_),
    .A3(\mod.Arithmetic.CN.I_in[30] ),
    .Z(_1313_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4643_ (.I(\mod.Arithmetic.CN.I_in[30] ),
    .Z(_1314_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4644_ (.A1(_1063_),
    .A2(_1178_),
    .B(_1314_),
    .ZN(_1315_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _4645_ (.A1(_1061_),
    .A2(_1313_),
    .A3(_1315_),
    .ZN(_1316_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _4646_ (.A1(_1312_),
    .A2(_1316_),
    .ZN(_1317_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _4647_ (.A1(_1174_),
    .A2(_1309_),
    .A3(_1317_),
    .Z(_1318_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _4648_ (.A1(_1306_),
    .A2(_1318_),
    .ZN(_1319_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4649_ (.A1(_1303_),
    .A2(_1319_),
    .Z(_1320_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4650_ (.A1(_1302_),
    .A2(_1320_),
    .Z(_1321_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _4651_ (.A1(_1297_),
    .A2(_1300_),
    .A3(_1321_),
    .ZN(_1322_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _4652_ (.A1(_1286_),
    .A2(_1322_),
    .ZN(_1323_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _4653_ (.A1(_1285_),
    .A2(_1323_),
    .ZN(_1324_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _4654_ (.A1(_1222_),
    .A2(_1256_),
    .Z(_1325_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _4655_ (.A1(_1222_),
    .A2(_1256_),
    .Z(_1326_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4656_ (.A1(_1219_),
    .A2(_1325_),
    .B(_1326_),
    .ZN(_1327_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4657_ (.A1(_1206_),
    .A2(_1212_),
    .ZN(_1328_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4658_ (.A1(_1208_),
    .A2(_1207_),
    .B1(_1328_),
    .B2(_1217_),
    .ZN(_1329_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4659_ (.I(\mod.Arithmetic.CN.I_in[37] ),
    .ZN(_1330_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _4660_ (.A1(_0651_),
    .A2(\mod.Arithmetic.CN.I_in[35] ),
    .A3(_1090_),
    .A4(_1330_),
    .ZN(_1331_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4661_ (.A1(_1090_),
    .A2(_1330_),
    .B(_1331_),
    .ZN(_1332_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4662_ (.A1(\mod.Arithmetic.CN.I_in[38] ),
    .A2(_1332_),
    .B(_1251_),
    .ZN(_1333_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4663_ (.A1(\mod.Arithmetic.CN.I_in[38] ),
    .A2(_1332_),
    .B(_1333_),
    .ZN(_1334_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4664_ (.A1(_1202_),
    .A2(\mod.Arithmetic.CN.I_in[45] ),
    .ZN(_1335_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4665_ (.A1(\mod.Arithmetic.CN.I_in[46] ),
    .A2(_1335_),
    .Z(_1336_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4666_ (.A1(_1251_),
    .A2(_1336_),
    .ZN(_1337_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4667_ (.I(\mod.Arithmetic.CN.I_in[45] ),
    .Z(_1338_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _4668_ (.A1(_1203_),
    .A2(_1338_),
    .A3(_0984_),
    .ZN(_1339_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4669_ (.A1(\mod.Arithmetic.CN.I_in[46] ),
    .A2(_1339_),
    .ZN(_1340_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4670_ (.A1(_1339_),
    .A2(_1337_),
    .B(_1340_),
    .ZN(_1341_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4671_ (.A1(_1338_),
    .A2(_1209_),
    .ZN(_1342_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _4672_ (.I0(_1337_),
    .I1(_1341_),
    .S(_1342_),
    .Z(_1343_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4673_ (.A1(_1334_),
    .A2(_1343_),
    .Z(_1344_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _4674_ (.A1(_1234_),
    .A2(_1344_),
    .ZN(_1345_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _4675_ (.A1(_1329_),
    .A2(_1345_),
    .ZN(_1346_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4676_ (.I(_1346_),
    .ZN(_1347_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4677_ (.A1(_1237_),
    .A2(_1254_),
    .ZN(_1348_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4678_ (.A1(_1236_),
    .A2(_1255_),
    .B(_1348_),
    .ZN(_1349_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _4679_ (.A1(_1224_),
    .A2(_1232_),
    .Z(_1350_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4680_ (.A1(_1227_),
    .A2(_1230_),
    .ZN(_1351_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _4681_ (.A1(_1225_),
    .A2(_0995_),
    .A3(_1231_),
    .B(_1351_),
    .ZN(_1352_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4682_ (.A1(\mod.Arithmetic.CN.I_in[61] ),
    .A2(_1135_),
    .ZN(_1353_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4683_ (.I(\mod.Arithmetic.CN.I_in[53] ),
    .ZN(_1354_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4684_ (.A1(\mod.Arithmetic.CN.I_in[52] ),
    .A2(_1354_),
    .ZN(_1355_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4685_ (.A1(\mod.Arithmetic.CN.I_in[54] ),
    .A2(_1355_),
    .Z(_1356_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _4686_ (.A1(_0636_),
    .A2(_1356_),
    .Z(_1357_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4687_ (.A1(_1353_),
    .A2(_1356_),
    .ZN(_1358_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4688_ (.A1(_1353_),
    .A2(_1357_),
    .B(_1358_),
    .ZN(_1359_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _4689_ (.A1(_1225_),
    .A2(_1354_),
    .A3(_0997_),
    .ZN(_1360_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4690_ (.A1(_1359_),
    .A2(_1360_),
    .Z(_1361_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4691_ (.A1(_1352_),
    .A2(_1361_),
    .Z(_1362_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4692_ (.A1(_1350_),
    .A2(_1362_),
    .Z(_1363_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _4693_ (.A1(_1240_),
    .A2(_1248_),
    .Z(_1364_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4694_ (.A1(_1249_),
    .A2(_1253_),
    .B(_1364_),
    .ZN(_1365_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4695_ (.I(\mod.Arithmetic.CN.I_in[62] ),
    .ZN(_1366_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4696_ (.A1(_1134_),
    .A2(_1250_),
    .B(_1366_),
    .ZN(_1367_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _4697_ (.A1(_1134_),
    .A2(_1250_),
    .A3(_1366_),
    .Z(_1368_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _4698_ (.A1(_0620_),
    .A2(_1367_),
    .A3(_1368_),
    .ZN(_1369_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _4699_ (.A1(_0891_),
    .A2(\mod.Arithmetic.CN.I_in[69] ),
    .Z(_1370_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4700_ (.A1(_1242_),
    .A2(_1246_),
    .ZN(_1371_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4701_ (.A1(_1370_),
    .A2(_1247_),
    .B(_1371_),
    .ZN(_1372_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4702_ (.A1(_0643_),
    .A2(\mod.Arithmetic.CN.I_in[70] ),
    .ZN(_1373_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _4703_ (.A1(\mod.Arithmetic.CN.I_in[67] ),
    .A2(_1245_),
    .B(_0634_),
    .C(\mod.Arithmetic.ACTI.x[4] ),
    .ZN(_1374_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _4704_ (.A1(_0641_),
    .A2(\mod.Arithmetic.ACTI.x[5] ),
    .A3(_1125_),
    .ZN(_1375_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4705_ (.A1(_0632_),
    .A2(\mod.Arithmetic.ACTI.x[6] ),
    .ZN(_1376_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4706_ (.A1(_1241_),
    .A2(_1376_),
    .Z(_1377_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4707_ (.A1(_1375_),
    .A2(_1377_),
    .Z(_1378_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4708_ (.A1(_1374_),
    .A2(_1378_),
    .Z(_1379_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4709_ (.A1(_1373_),
    .A2(_1379_),
    .Z(_1380_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4710_ (.A1(_1372_),
    .A2(_1380_),
    .Z(_1381_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _4711_ (.A1(_1369_),
    .A2(_1381_),
    .ZN(_1382_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4712_ (.A1(_1365_),
    .A2(_1382_),
    .Z(_1383_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _4713_ (.A1(_1363_),
    .A2(_1383_),
    .ZN(_1384_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _4714_ (.A1(_1349_),
    .A2(_1384_),
    .ZN(_1385_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4715_ (.A1(_1347_),
    .A2(_1385_),
    .Z(_1386_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _4716_ (.A1(_1324_),
    .A2(_1327_),
    .A3(_1386_),
    .ZN(_1387_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _4717_ (.A1(_1279_),
    .A2(_1282_),
    .A3(_1387_),
    .ZN(_1388_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4718_ (.A1(_1276_),
    .A2(_1388_),
    .Z(_1389_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _4719_ (.A1(_1273_),
    .A2(_1389_),
    .ZN(_1390_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _4720_ (.A1(_1272_),
    .A2(_1390_),
    .ZN(_1391_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _4721_ (.A1(_1269_),
    .A2(_1391_),
    .Z(_1392_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4722_ (.A1(_1269_),
    .A2(_1391_),
    .ZN(_1393_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _4723_ (.A1(_1031_),
    .A2(_1392_),
    .A3(_1393_),
    .ZN(_1394_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4724_ (.A1(_0789_),
    .A2(_1266_),
    .B(_1268_),
    .C(_1394_),
    .ZN(\mod.P3.Res[6] ));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _4725_ (.A1(_1272_),
    .A2(_1390_),
    .Z(_1395_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4726_ (.A1(_1276_),
    .A2(_1388_),
    .B1(_1389_),
    .B2(_1273_),
    .ZN(_1396_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4727_ (.A1(_1282_),
    .A2(_1387_),
    .ZN(_1397_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4728_ (.A1(_1282_),
    .A2(_1387_),
    .ZN(_1398_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4729_ (.A1(_1279_),
    .A2(_1397_),
    .B(_1398_),
    .ZN(_1399_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4730_ (.I(_1349_),
    .ZN(_1400_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4731_ (.A1(_1347_),
    .A2(_1385_),
    .ZN(_1401_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4732_ (.A1(_1400_),
    .A2(_1384_),
    .B(_1401_),
    .ZN(_1402_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4733_ (.A1(\mod.Arithmetic.CN.I_in[61] ),
    .A2(_1366_),
    .ZN(_1403_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4734_ (.A1(\mod.Arithmetic.CN.I_in[63] ),
    .A2(_1403_),
    .Z(_1404_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4735_ (.A1(_0625_),
    .A2(_1404_),
    .ZN(_1405_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _4736_ (.A1(_1293_),
    .A2(_1402_),
    .A3(_1405_),
    .Z(_1406_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4737_ (.A1(_1350_),
    .A2(_1362_),
    .ZN(_1407_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _4738_ (.A1(_1338_),
    .A2(_1209_),
    .A3(_1337_),
    .ZN(_1408_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4739_ (.A1(_1334_),
    .A2(_1343_),
    .B(_1408_),
    .ZN(_1409_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4740_ (.A1(_1407_),
    .A2(_1409_),
    .Z(_1410_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4741_ (.I(_1338_),
    .ZN(_1411_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4742_ (.A1(_1411_),
    .A2(\mod.Arithmetic.CN.I_in[46] ),
    .ZN(_1412_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _4743_ (.A1(\mod.Arithmetic.CN.I_in[47] ),
    .A2(_1412_),
    .ZN(_1413_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4744_ (.A1(_0622_),
    .A2(_1413_),
    .ZN(_1414_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4745_ (.A1(_0622_),
    .A2(\mod.Arithmetic.CN.I_in[71] ),
    .ZN(_1415_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4746_ (.A1(\mod.Arithmetic.CN.I_in[69] ),
    .A2(_1376_),
    .ZN(_1416_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _4747_ (.I0(_1373_),
    .I1(\mod.Arithmetic.CN.I_in[70] ),
    .S(_1416_),
    .Z(_1417_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _4748_ (.A1(_1414_),
    .A2(_1415_),
    .A3(_1417_),
    .Z(_1418_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _4749_ (.A1(_0623_),
    .A2(\mod.Arithmetic.CN.I_in[70] ),
    .A3(_1379_),
    .ZN(_1419_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4750_ (.A1(_1374_),
    .A2(_1378_),
    .B(_1419_),
    .ZN(_1420_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _4751_ (.A1(_1203_),
    .A2(\mod.Arithmetic.CN.I_in[46] ),
    .A3(_1208_),
    .B(_1340_),
    .ZN(_1421_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4752_ (.I(_0623_),
    .Z(_1422_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4753_ (.I(\mod.Arithmetic.CN.I_in[38] ),
    .ZN(_1423_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4754_ (.A1(_1185_),
    .A2(_1423_),
    .ZN(_1424_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _4755_ (.A1(\mod.Arithmetic.CN.I_in[37] ),
    .A2(_1423_),
    .B1(_1213_),
    .B2(_1424_),
    .ZN(_1425_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4756_ (.A1(\mod.Arithmetic.CN.I_in[39] ),
    .A2(_1425_),
    .Z(_1426_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4757_ (.A1(_1422_),
    .A2(_1426_),
    .ZN(_1427_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4758_ (.A1(_1421_),
    .A2(_1427_),
    .Z(_1428_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _4759_ (.A1(_1418_),
    .A2(_1420_),
    .A3(_1428_),
    .Z(_1429_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4760_ (.A1(_1286_),
    .A2(_1322_),
    .ZN(_1430_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4761_ (.A1(_1285_),
    .A2(_1323_),
    .B(_1430_),
    .ZN(_1431_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _4762_ (.A1(_1410_),
    .A2(_1429_),
    .A3(_1431_),
    .Z(_1432_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _4763_ (.A1(_1251_),
    .A2(_1354_),
    .A3(\mod.Arithmetic.CN.I_in[54] ),
    .ZN(_1433_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4764_ (.A1(_1352_),
    .A2(_1361_),
    .B1(_1433_),
    .B2(_1225_),
    .ZN(_1434_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4765_ (.A1(_1359_),
    .A2(_1360_),
    .B(_1434_),
    .C(_1358_),
    .ZN(_1435_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4766_ (.A1(_1422_),
    .A2(\mod.Arithmetic.ACTI.x[7] ),
    .ZN(_1436_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _4767_ (.A1(\mod.Arithmetic.CN.I_in[68] ),
    .A2(_1377_),
    .B(_1422_),
    .C(\mod.Arithmetic.ACTI.x[5] ),
    .ZN(_1437_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _4768_ (.I0(\mod.Arithmetic.ACTI.x[7] ),
    .I1(_1436_),
    .S(_1437_),
    .Z(_1438_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _4769_ (.A1(_0624_),
    .A2(_1134_),
    .A3(\mod.Arithmetic.CN.I_in[61] ),
    .A4(_1366_),
    .ZN(_1439_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4770_ (.A1(_0624_),
    .A2(_1439_),
    .ZN(_1440_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4771_ (.A1(_1354_),
    .A2(\mod.Arithmetic.CN.I_in[54] ),
    .ZN(_1441_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4772_ (.A1(\mod.Arithmetic.CN.I_in[55] ),
    .A2(_1441_),
    .Z(_1442_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _4773_ (.I0(_1440_),
    .I1(_1439_),
    .S(_1442_),
    .Z(_1443_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _4774_ (.A1(_1435_),
    .A2(_1438_),
    .A3(_1443_),
    .Z(_1444_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4775_ (.A1(_1300_),
    .A2(_1321_),
    .ZN(_1445_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4776_ (.A1(_1300_),
    .A2(_1321_),
    .ZN(_1446_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4777_ (.A1(_1297_),
    .A2(_1445_),
    .B(_1446_),
    .ZN(_1447_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4778_ (.A1(_1309_),
    .A2(_1317_),
    .ZN(_1448_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _4779_ (.A1(_1306_),
    .A2(_1318_),
    .Z(_1449_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4780_ (.A1(_1309_),
    .A2(_1317_),
    .ZN(_1450_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _4781_ (.A1(_1174_),
    .A2(_1448_),
    .B(_1449_),
    .C(_1450_),
    .ZN(_1451_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4782_ (.A1(_1447_),
    .A2(_1451_),
    .Z(_1452_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _4783_ (.A1(_0743_),
    .A2(_1190_),
    .A3(_1188_),
    .ZN(_1453_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4784_ (.A1(_0743_),
    .A2(_1294_),
    .B(_1453_),
    .ZN(_1454_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4785_ (.A1(_1288_),
    .A2(_0735_),
    .ZN(_1455_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4786_ (.A1(\mod.Arithmetic.CN.I_in[15] ),
    .A2(_1455_),
    .Z(_1456_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4787_ (.A1(_0624_),
    .A2(_1456_),
    .ZN(_1457_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4788_ (.A1(_1234_),
    .A2(_1344_),
    .ZN(_1458_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4789_ (.A1(_1329_),
    .A2(_1345_),
    .B(_1458_),
    .ZN(_1459_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4790_ (.A1(_1307_),
    .A2(_1314_),
    .ZN(_1460_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4791_ (.A1(\mod.Arithmetic.CN.I_in[23] ),
    .A2(\mod.Arithmetic.CN.I_in[31] ),
    .Z(_1461_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _4792_ (.A1(_0696_),
    .A2(_1460_),
    .A3(_1461_),
    .Z(_1462_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4793_ (.A1(_1422_),
    .A2(_1462_),
    .ZN(_1463_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _4794_ (.A1(_1423_),
    .A2(_1331_),
    .Z(_1464_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4795_ (.A1(_1303_),
    .A2(_1319_),
    .ZN(_1465_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4796_ (.A1(_1302_),
    .A2(_1320_),
    .B(_1465_),
    .ZN(_1466_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4797_ (.A1(_1312_),
    .A2(_1316_),
    .ZN(_1467_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4798_ (.A1(_1314_),
    .A2(_1176_),
    .B(_1310_),
    .C(_1467_),
    .ZN(_1468_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _4799_ (.A1(_1314_),
    .A2(_1176_),
    .A3(_1310_),
    .B(_1468_),
    .ZN(_1469_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _4800_ (.A1(_1464_),
    .A2(_1466_),
    .A3(_1469_),
    .ZN(_1470_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _4801_ (.A1(_1459_),
    .A2(_1463_),
    .A3(_1470_),
    .Z(_1471_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _4802_ (.A1(_1454_),
    .A2(_1457_),
    .A3(_1471_),
    .Z(_1472_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _4803_ (.A1(_1444_),
    .A2(_1452_),
    .A3(_1472_),
    .Z(_1473_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _4804_ (.A1(_1406_),
    .A2(_1432_),
    .A3(_1473_),
    .Z(_1474_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4805_ (.A1(_1327_),
    .A2(_1386_),
    .ZN(_1475_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4806_ (.A1(_1327_),
    .A2(_1386_),
    .ZN(_1476_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4807_ (.A1(_1324_),
    .A2(_1475_),
    .B(_1476_),
    .ZN(_1477_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _4808_ (.A1(_0625_),
    .A2(_1367_),
    .A3(_1368_),
    .A4(_1381_),
    .ZN(_1478_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4809_ (.A1(_1372_),
    .A2(_1380_),
    .B(_1478_),
    .ZN(_1479_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _4810_ (.A1(_1365_),
    .A2(_1382_),
    .Z(_1480_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4811_ (.A1(_1363_),
    .A2(_1383_),
    .B(_1480_),
    .ZN(_1481_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _4812_ (.A1(_1477_),
    .A2(_1479_),
    .A3(_1481_),
    .Z(_1482_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _4813_ (.A1(_1399_),
    .A2(_1474_),
    .A3(_1482_),
    .Z(_1483_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4814_ (.A1(_1396_),
    .A2(_1483_),
    .Z(_1484_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _4815_ (.A1(_1395_),
    .A2(_1392_),
    .A3(_1484_),
    .Z(_1485_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4816_ (.A1(_1395_),
    .A2(_1392_),
    .B(_1484_),
    .ZN(_1486_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4817_ (.A1(_0797_),
    .A2(_0672_),
    .ZN(_1487_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_1 _4818_ (.A1(_0673_),
    .A2(_0674_),
    .A3(\mod.Arithmetic.I_out[79] ),
    .A4(_0675_),
    .ZN(_1488_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _4819_ (.A1(_1267_),
    .A2(_1485_),
    .A3(_1486_),
    .B1(_1487_),
    .B2(_1488_),
    .ZN(\mod.P3.Res[7] ));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4820_ (.I(\mod.Data_Mem.F_M.src[8] ),
    .Z(_1489_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4821_ (.I(_1489_),
    .Z(_1490_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4822_ (.I(_1490_),
    .Z(_1491_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4823_ (.I(\mod.Data_Mem.F_M.src[1] ),
    .ZN(_1492_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4824_ (.I(_1492_),
    .Z(_1493_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4825_ (.I(\mod.Data_Mem.F_M.src[2] ),
    .Z(_1494_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4826_ (.I(\mod.Data_Mem.F_M.src[4] ),
    .Z(_1495_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4827_ (.A1(_1494_),
    .A2(_1495_),
    .ZN(_1496_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4828_ (.A1(_1493_),
    .A2(_1496_),
    .ZN(_1497_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4829_ (.I(_1497_),
    .Z(_1498_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4830_ (.I(_1495_),
    .Z(_1499_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4831_ (.I(\mod.Data_Mem.F_M.src[2] ),
    .ZN(_1500_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4832_ (.I(_1500_),
    .Z(_1501_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4833_ (.I(\mod.Data_Mem.F_M.src[0] ),
    .Z(_1502_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4834_ (.I(\mod.Data_Mem.F_M.src[1] ),
    .Z(_1503_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4835_ (.A1(_1502_),
    .A2(_1503_),
    .ZN(_1504_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4836_ (.A1(_1501_),
    .A2(_1504_),
    .ZN(_1505_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4837_ (.A1(_1499_),
    .A2(_1505_),
    .ZN(_1506_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4838_ (.I(_1506_),
    .Z(_1507_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4839_ (.I(_1507_),
    .Z(_1508_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4840_ (.I(_1502_),
    .Z(_1509_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _4841_ (.I(_1509_),
    .Z(_1510_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _4842_ (.I0(\mod.Data_Mem.F_M.MRAM[21][0] ),
    .I1(\mod.Data_Mem.F_M.MRAM[20][0] ),
    .S(_1510_),
    .Z(_1511_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4843_ (.I(_1502_),
    .Z(_1512_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4844_ (.I(_1512_),
    .Z(_1513_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4845_ (.I(_1513_),
    .Z(_1514_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _4846_ (.I(_1514_),
    .Z(_1515_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _4847_ (.I0(\mod.Data_Mem.F_M.MRAM[19][0] ),
    .I1(\mod.Data_Mem.F_M.MRAM[18][0] ),
    .S(_1515_),
    .Z(_1516_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4848_ (.I(_1512_),
    .Z(_1517_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4849_ (.I(_1517_),
    .Z(_1518_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4850_ (.I(_1518_),
    .Z(_1519_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _4851_ (.I0(\mod.Data_Mem.F_M.MRAM[17][0] ),
    .I1(\mod.Data_Mem.F_M.MRAM[16][0] ),
    .S(_1519_),
    .Z(_1520_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4852_ (.I(\mod.Data_Mem.F_M.src[0] ),
    .ZN(_1521_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4853_ (.I(_1521_),
    .Z(_1522_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4854_ (.A1(_1522_),
    .A2(_1492_),
    .ZN(_1523_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4855_ (.A1(_1504_),
    .A2(_1523_),
    .ZN(_1524_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4856_ (.I(_1524_),
    .Z(_1525_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4857_ (.I(_1525_),
    .Z(_1526_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _4858_ (.I(_1526_),
    .Z(_1527_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4859_ (.A1(_1521_),
    .A2(_1492_),
    .ZN(_1528_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4860_ (.A1(_1501_),
    .A2(_1528_),
    .ZN(_1529_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4861_ (.I(_1529_),
    .Z(_1530_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4862_ (.I(_1530_),
    .Z(_1531_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _4863_ (.I0(\mod.Data_Mem.F_M.MRAM[22][0] ),
    .I1(_1511_),
    .I2(_1516_),
    .I3(_1520_),
    .S0(_1527_),
    .S1(_1531_),
    .Z(_1532_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4864_ (.I(_1496_),
    .Z(_1533_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4865_ (.I(\mod.Data_Mem.F_M.src[4] ),
    .ZN(_1534_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4866_ (.I(_1534_),
    .Z(_1535_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4867_ (.I(_1535_),
    .Z(_1536_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4868_ (.I(_1528_),
    .Z(_1537_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4869_ (.I(_1537_),
    .Z(_1538_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4870_ (.I(_1538_),
    .Z(_1539_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _4871_ (.I0(\mod.Data_Mem.F_M.MRAM[5][0] ),
    .I1(\mod.Data_Mem.F_M.MRAM[4][0] ),
    .S(_1514_),
    .Z(_1540_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4872_ (.A1(\mod.Data_Mem.F_M.src[0] ),
    .A2(_1503_),
    .ZN(_1541_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4873_ (.I(_1541_),
    .Z(_1542_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4874_ (.I(_1542_),
    .Z(_1543_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _4875_ (.I0(\mod.Data_Mem.F_M.MRAM[6][0] ),
    .I1(_1540_),
    .S(_1543_),
    .Z(_1544_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _4876_ (.A1(\mod.Data_Mem.F_M.MRAM[3][0] ),
    .A2(_1539_),
    .B1(_1531_),
    .B2(_1544_),
    .ZN(_1545_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4877_ (.A1(_1536_),
    .A2(_1545_),
    .ZN(_1546_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4878_ (.A1(_1508_),
    .A2(_1532_),
    .B(_1533_),
    .C(_1546_),
    .ZN(_1547_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4879_ (.I(_1494_),
    .Z(_1548_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4880_ (.I(_1504_),
    .Z(_1549_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4881_ (.A1(_1548_),
    .A2(_1549_),
    .ZN(_1550_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4882_ (.I(_1550_),
    .Z(_1551_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4883_ (.I(_1551_),
    .Z(_1552_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4884_ (.I(_1534_),
    .Z(_1553_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4885_ (.I(\mod.Data_Mem.F_M.src[2] ),
    .Z(_1554_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4886_ (.A1(_1554_),
    .A2(_1537_),
    .ZN(_1555_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4887_ (.A1(_1553_),
    .A2(_1555_),
    .ZN(_1556_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4888_ (.I(_1556_),
    .Z(_1557_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4889_ (.I(_1557_),
    .Z(_1558_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _4890_ (.A1(\mod.Data_Mem.F_M.MRAM[15][0] ),
    .A2(_1536_),
    .B1(\mod.Data_Mem.F_M.MRAM[31][0] ),
    .B2(_1558_),
    .C(_1551_),
    .ZN(_1559_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4891_ (.A1(_1547_),
    .A2(_1552_),
    .B(_1559_),
    .ZN(_1560_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4892_ (.A1(_1554_),
    .A2(_1504_),
    .ZN(_1561_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4893_ (.I(_1561_),
    .Z(_1562_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4894_ (.I(_1562_),
    .Z(_1563_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4895_ (.I(_1525_),
    .Z(_1564_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4896_ (.I(_1564_),
    .Z(_1565_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4897_ (.I(_1565_),
    .Z(_1566_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4898_ (.I(_1513_),
    .Z(_1567_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _4899_ (.I(_1567_),
    .Z(_1568_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _4900_ (.I0(\mod.Data_Mem.F_M.MRAM[773][0] ),
    .I1(\mod.Data_Mem.F_M.MRAM[772][0] ),
    .S(_1568_),
    .Z(_1569_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4901_ (.A1(_1566_),
    .A2(_1569_),
    .ZN(_1570_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4902_ (.A1(_1528_),
    .A2(_1541_),
    .ZN(_1571_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4903_ (.I(_1571_),
    .Z(_1572_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4904_ (.I(_1572_),
    .Z(_1573_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4905_ (.I(_1573_),
    .Z(_1574_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4906_ (.I(_1574_),
    .Z(_1575_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4907_ (.A1(\mod.Data_Mem.F_M.MRAM[774][0] ),
    .A2(_1575_),
    .ZN(_1576_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _4908_ (.A1(_1563_),
    .A2(_1570_),
    .A3(_1576_),
    .ZN(_1577_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4909_ (.I(_1502_),
    .Z(_1578_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4910_ (.I(_1578_),
    .Z(_1579_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4911_ (.I(_1579_),
    .Z(_1580_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4912_ (.I(_1580_),
    .Z(_1581_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _4913_ (.I0(\mod.Data_Mem.F_M.MRAM[771][0] ),
    .I1(\mod.Data_Mem.F_M.MRAM[770][0] ),
    .S(_1581_),
    .Z(_1582_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4914_ (.A1(_1575_),
    .A2(_1582_),
    .ZN(_1583_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4915_ (.I(_1564_),
    .Z(_1584_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4916_ (.I(_1584_),
    .Z(_1585_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4917_ (.I(_1578_),
    .Z(_1586_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4918_ (.I(_1586_),
    .Z(_1587_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4919_ (.I(_1587_),
    .Z(_1588_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _4920_ (.I0(\mod.Data_Mem.F_M.MRAM[769][0] ),
    .I1(\mod.Data_Mem.F_M.MRAM[768][0] ),
    .S(_1588_),
    .Z(_1589_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4921_ (.I(_1561_),
    .Z(_1590_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4922_ (.A1(_1585_),
    .A2(_1589_),
    .B(_1590_),
    .ZN(_1591_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4923_ (.A1(_1583_),
    .A2(_1591_),
    .B(_1558_),
    .ZN(_1592_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4924_ (.I(_1512_),
    .Z(_1593_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4925_ (.I(_1593_),
    .Z(_1594_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4926_ (.I(_1492_),
    .Z(_1595_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4927_ (.A1(_1595_),
    .A2(_1494_),
    .ZN(_1596_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4928_ (.A1(_1594_),
    .A2(_1596_),
    .ZN(_1597_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4929_ (.I(_1597_),
    .Z(_1598_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4930_ (.I(_1598_),
    .Z(_1599_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4931_ (.I(_1523_),
    .Z(_1600_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4932_ (.I(_1600_),
    .Z(_1601_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4933_ (.I(_1525_),
    .Z(_1602_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4934_ (.I(_1602_),
    .Z(_1603_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _4935_ (.I0(\mod.Data_Mem.F_M.MRAM[789][0] ),
    .I1(\mod.Data_Mem.F_M.MRAM[788][0] ),
    .S(_1568_),
    .Z(_1604_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4936_ (.A1(\mod.Data_Mem.F_M.MRAM[790][0] ),
    .A2(_1601_),
    .B1(_1603_),
    .B2(_1604_),
    .ZN(_1605_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4937_ (.I(_1572_),
    .Z(_1606_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4938_ (.I(_1606_),
    .Z(_1607_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4939_ (.I(_1607_),
    .Z(_1608_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4940_ (.I(_1509_),
    .Z(_1609_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _4941_ (.I0(\mod.Data_Mem.F_M.MRAM[787][0] ),
    .I1(\mod.Data_Mem.F_M.MRAM[786][0] ),
    .S(_1609_),
    .Z(_1610_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4942_ (.A1(_1608_),
    .A2(_1610_),
    .ZN(_1611_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4943_ (.I(_1567_),
    .Z(_1612_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _4944_ (.I0(\mod.Data_Mem.F_M.MRAM[785][0] ),
    .I1(\mod.Data_Mem.F_M.MRAM[784][0] ),
    .S(_1612_),
    .Z(_1613_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4945_ (.I(_1561_),
    .Z(_1614_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4946_ (.A1(_1603_),
    .A2(_1613_),
    .B(_1614_),
    .ZN(_1615_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4947_ (.I(_1506_),
    .Z(_1616_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _4948_ (.A1(_1563_),
    .A2(_1605_),
    .B1(_1611_),
    .B2(_1615_),
    .C(_1616_),
    .ZN(_1617_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _4949_ (.A1(_1577_),
    .A2(_1592_),
    .B(_1599_),
    .C(_1617_),
    .ZN(_1618_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4950_ (.I(_1499_),
    .Z(_1619_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4951_ (.I(_1619_),
    .Z(_1620_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4952_ (.I(_1507_),
    .Z(_1621_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4953_ (.I(_1550_),
    .Z(_1622_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _4954_ (.A1(_1620_),
    .A2(\mod.Data_Mem.F_M.MRAM[799][0] ),
    .B1(_1621_),
    .B2(\mod.Data_Mem.F_M.MRAM[783][0] ),
    .C(_1622_),
    .ZN(_1623_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4955_ (.A1(_1618_),
    .A2(_1623_),
    .ZN(_1624_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4956_ (.I(_1489_),
    .Z(_1625_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4957_ (.A1(_1501_),
    .A2(_1553_),
    .ZN(_1626_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4958_ (.I(_1626_),
    .Z(_1627_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4959_ (.A1(_1539_),
    .A2(_1627_),
    .ZN(_1628_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4960_ (.A1(_1625_),
    .A2(_1628_),
    .ZN(_1629_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _4961_ (.A1(_1491_),
    .A2(_1498_),
    .A3(_1560_),
    .B1(_1624_),
    .B2(_1629_),
    .ZN(_1630_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4962_ (.I(_1630_),
    .ZN(_0000_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4963_ (.I(_1628_),
    .Z(_1631_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4964_ (.I(\mod.Data_Mem.F_M.MRAM[31][1] ),
    .Z(_1632_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4965_ (.I(_1616_),
    .Z(_1633_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4966_ (.A1(_1620_),
    .A2(_1632_),
    .B1(_1633_),
    .B2(\mod.Data_Mem.F_M.MRAM[15][1] ),
    .ZN(_1634_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4967_ (.I(_1584_),
    .Z(_1635_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4968_ (.I(_1594_),
    .Z(_1636_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _4969_ (.I0(\mod.Data_Mem.F_M.MRAM[5][1] ),
    .I1(\mod.Data_Mem.F_M.MRAM[4][1] ),
    .S(_1636_),
    .Z(_1637_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4970_ (.A1(_1635_),
    .A2(_1637_),
    .ZN(_1638_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4971_ (.I(_1600_),
    .Z(_1639_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4972_ (.I(_1639_),
    .Z(_1640_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4973_ (.I(_1529_),
    .Z(_1641_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4974_ (.I(_1641_),
    .Z(_1642_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4975_ (.A1(\mod.Data_Mem.F_M.MRAM[6][1] ),
    .A2(_1640_),
    .B(_1642_),
    .ZN(_1643_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4976_ (.I(_1606_),
    .Z(_1644_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4977_ (.I(_1644_),
    .Z(_1645_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4978_ (.I(_1593_),
    .Z(_1646_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4979_ (.I(_1646_),
    .Z(_1647_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _4980_ (.I0(\mod.Data_Mem.F_M.MRAM[3][1] ),
    .I1(\mod.Data_Mem.F_M.MRAM[2][1] ),
    .S(_1647_),
    .Z(_1648_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _4981_ (.I0(\mod.Data_Mem.F_M.MRAM[1][1] ),
    .I1(\mod.Data_Mem.F_M.MRAM[0][1] ),
    .S(_1509_),
    .Z(_1649_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _4982_ (.A1(_1565_),
    .A2(_1649_),
    .Z(_1650_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4983_ (.I(_1561_),
    .Z(_1651_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _4984_ (.A1(_1645_),
    .A2(_1648_),
    .B(_1650_),
    .C(_1651_),
    .ZN(_1652_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4985_ (.I(_1556_),
    .Z(_1653_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _4986_ (.A1(_1638_),
    .A2(_1643_),
    .B(_1652_),
    .C(_1653_),
    .ZN(_1654_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4987_ (.I(_1584_),
    .Z(_1655_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _4988_ (.I0(\mod.Data_Mem.F_M.MRAM[17][1] ),
    .I1(\mod.Data_Mem.F_M.MRAM[16][1] ),
    .S(_1519_),
    .Z(_1656_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4989_ (.A1(_1655_),
    .A2(_1656_),
    .ZN(_1657_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4990_ (.I(_1646_),
    .Z(_1658_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _4991_ (.I0(\mod.Data_Mem.F_M.MRAM[19][1] ),
    .I1(\mod.Data_Mem.F_M.MRAM[18][1] ),
    .S(_1658_),
    .Z(_1659_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4992_ (.A1(_1608_),
    .A2(_1659_),
    .B(_1614_),
    .ZN(_1660_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4993_ (.I(_1639_),
    .Z(_1661_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4994_ (.A1(\mod.Data_Mem.F_M.MRAM[22][1] ),
    .A2(_1661_),
    .B(_1531_),
    .ZN(_1662_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4995_ (.I(_1525_),
    .Z(_1663_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4996_ (.I(_1663_),
    .Z(_1664_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _4997_ (.I0(\mod.Data_Mem.F_M.MRAM[21][1] ),
    .I1(\mod.Data_Mem.F_M.MRAM[20][1] ),
    .S(_1636_),
    .Z(_1665_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4998_ (.A1(_1664_),
    .A2(_1665_),
    .ZN(_1666_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _4999_ (.A1(_1657_),
    .A2(_1660_),
    .B1(_1662_),
    .B2(_1666_),
    .C(_1616_),
    .ZN(_1667_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5000_ (.A1(_1654_),
    .A2(_1667_),
    .B(_1622_),
    .ZN(_1668_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5001_ (.I(\mod.Data_Mem.F_M.src[8] ),
    .ZN(_1669_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5002_ (.I(_1669_),
    .Z(_1670_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _5003_ (.A1(_1552_),
    .A2(_1634_),
    .B(_1668_),
    .C(_1670_),
    .ZN(_1671_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5004_ (.I(_1598_),
    .Z(_1672_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5005_ (.I(_1672_),
    .Z(_1673_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5006_ (.I(_1598_),
    .Z(_1674_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5007_ (.I(_1514_),
    .Z(_1675_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5008_ (.I(_1593_),
    .Z(_1676_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5009_ (.I(_1676_),
    .Z(_1677_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5010_ (.I(\mod.Data_Mem.F_M.MRAM[784][1] ),
    .ZN(_1678_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5011_ (.A1(_1677_),
    .A2(_1678_),
    .ZN(_1679_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5012_ (.A1(_1675_),
    .A2(\mod.Data_Mem.F_M.MRAM[785][1] ),
    .B(_1679_),
    .ZN(_1680_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5013_ (.I(_1676_),
    .Z(_1681_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5014_ (.I(\mod.Data_Mem.F_M.MRAM[786][1] ),
    .ZN(_1682_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5015_ (.A1(_1681_),
    .A2(_1682_),
    .ZN(_1683_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5016_ (.A1(_1675_),
    .A2(\mod.Data_Mem.F_M.MRAM[787][1] ),
    .B(_1683_),
    .ZN(_1684_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5017_ (.I(_1518_),
    .Z(_1685_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5018_ (.I(_1594_),
    .Z(_1686_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5019_ (.I(\mod.Data_Mem.F_M.MRAM[788][1] ),
    .ZN(_1687_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5020_ (.A1(_1686_),
    .A2(_1687_),
    .ZN(_1688_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5021_ (.A1(_1685_),
    .A2(\mod.Data_Mem.F_M.MRAM[789][1] ),
    .B(_1688_),
    .ZN(_1689_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5022_ (.I(_1522_),
    .Z(_1690_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5023_ (.I(_1690_),
    .Z(_1691_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5024_ (.I(_1579_),
    .Z(_1692_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _5025_ (.A1(_1692_),
    .A2(\mod.Data_Mem.F_M.MRAM[790][1] ),
    .Z(_1693_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5026_ (.A1(_1691_),
    .A2(\mod.Data_Mem.F_M.MRAM[791][1] ),
    .B(_1693_),
    .ZN(_1694_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5027_ (.I(_1571_),
    .Z(_1695_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _5028_ (.I0(_1680_),
    .I1(_1684_),
    .I2(_1689_),
    .I3(_1694_),
    .S0(_1695_),
    .S1(_1651_),
    .Z(_1696_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5029_ (.A1(_1674_),
    .A2(_1696_),
    .B(_1558_),
    .ZN(_1697_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5030_ (.A1(\mod.Data_Mem.F_M.MRAM[799][1] ),
    .A2(_1673_),
    .B(_1697_),
    .ZN(_1698_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5031_ (.I(_1672_),
    .Z(_1699_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5032_ (.I(_1562_),
    .Z(_1700_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _5033_ (.I(_1676_),
    .Z(_1701_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5034_ (.I0(\mod.Data_Mem.F_M.MRAM[773][1] ),
    .I1(\mod.Data_Mem.F_M.MRAM[772][1] ),
    .S(_1701_),
    .Z(_1702_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5035_ (.I0(\mod.Data_Mem.F_M.MRAM[775][1] ),
    .I1(\mod.Data_Mem.F_M.MRAM[774][1] ),
    .S(_1692_),
    .Z(_1703_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5036_ (.I(_1573_),
    .Z(_1704_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5037_ (.I0(_1702_),
    .I1(_1703_),
    .S(_1704_),
    .Z(_1705_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5038_ (.I(_1644_),
    .Z(_1706_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5039_ (.I(_1567_),
    .Z(_1707_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5040_ (.I(_1512_),
    .Z(_1708_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5041_ (.I(\mod.Data_Mem.F_M.MRAM[770][1] ),
    .ZN(_1709_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5042_ (.A1(_1708_),
    .A2(_1709_),
    .ZN(_1710_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5043_ (.A1(_1707_),
    .A2(\mod.Data_Mem.F_M.MRAM[771][1] ),
    .B(_1710_),
    .ZN(_1711_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5044_ (.A1(_1706_),
    .A2(_1711_),
    .ZN(_1712_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5045_ (.I(_1526_),
    .Z(_1713_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5046_ (.I(_1578_),
    .Z(_1714_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5047_ (.I(_1646_),
    .Z(_1715_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5048_ (.I(\mod.Data_Mem.F_M.MRAM[768][1] ),
    .ZN(_1716_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5049_ (.A1(_1715_),
    .A2(_1716_),
    .ZN(_1717_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5050_ (.A1(_1714_),
    .A2(\mod.Data_Mem.F_M.MRAM[769][1] ),
    .B(_1717_),
    .ZN(_1718_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5051_ (.A1(_1713_),
    .A2(_1718_),
    .B(_1651_),
    .ZN(_1719_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5052_ (.A1(_1700_),
    .A2(_1705_),
    .B1(_1712_),
    .B2(_1719_),
    .ZN(_1720_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5053_ (.I(_1507_),
    .Z(_1721_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5054_ (.A1(_1674_),
    .A2(_1720_),
    .B(_1721_),
    .ZN(_1722_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5055_ (.A1(\mod.Data_Mem.F_M.MRAM[783][1] ),
    .A2(_1699_),
    .B(_1722_),
    .ZN(_1723_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5056_ (.I(\mod.Data_Mem.F_M.src[8] ),
    .Z(_1724_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5057_ (.I(_1724_),
    .Z(_1725_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5058_ (.I(_1725_),
    .Z(_1726_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5059_ (.A1(_1698_),
    .A2(_1723_),
    .B(_1726_),
    .ZN(_1727_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _5060_ (.A1(_1631_),
    .A2(_1671_),
    .A3(_1727_),
    .ZN(_1728_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5061_ (.I(_1728_),
    .ZN(_0001_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5062_ (.I(_1537_),
    .Z(_1729_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5063_ (.I(_1602_),
    .Z(_1730_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5064_ (.I0(\mod.Data_Mem.F_M.MRAM[5][2] ),
    .I1(\mod.Data_Mem.F_M.MRAM[4][2] ),
    .S(_1636_),
    .Z(_1731_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5065_ (.A1(_1730_),
    .A2(_1731_),
    .ZN(_1732_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5066_ (.A1(\mod.Data_Mem.F_M.MRAM[6][2] ),
    .A2(_1601_),
    .B(_1641_),
    .ZN(_1733_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5067_ (.I(_1526_),
    .Z(_1734_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5068_ (.I0(\mod.Data_Mem.F_M.MRAM[1][2] ),
    .I1(\mod.Data_Mem.F_M.MRAM[0][2] ),
    .S(_1658_),
    .Z(_1735_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5069_ (.A1(_1734_),
    .A2(_1735_),
    .ZN(_1736_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5070_ (.I(_1606_),
    .Z(_1737_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _5071_ (.I(_1737_),
    .Z(_1738_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5072_ (.I0(\mod.Data_Mem.F_M.MRAM[3][2] ),
    .I1(\mod.Data_Mem.F_M.MRAM[2][2] ),
    .S(_1647_),
    .Z(_1739_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5073_ (.A1(_1738_),
    .A2(_1739_),
    .B(_1562_),
    .ZN(_1740_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5074_ (.A1(_1732_),
    .A2(_1733_),
    .B1(_1736_),
    .B2(_1740_),
    .ZN(_1741_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5075_ (.I(_1524_),
    .Z(_1742_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5076_ (.I0(\mod.Data_Mem.F_M.MRAM[17][2] ),
    .I1(\mod.Data_Mem.F_M.MRAM[16][2] ),
    .S(_1519_),
    .Z(_1743_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5077_ (.A1(_1742_),
    .A2(_1743_),
    .ZN(_1744_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5078_ (.I(_1572_),
    .Z(_1745_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _5079_ (.I(_1518_),
    .Z(_1746_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5080_ (.I0(\mod.Data_Mem.F_M.MRAM[19][2] ),
    .I1(\mod.Data_Mem.F_M.MRAM[18][2] ),
    .S(_1746_),
    .Z(_1747_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5081_ (.A1(_1745_),
    .A2(_1747_),
    .B(_1562_),
    .ZN(_1748_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _5082_ (.I(_1600_),
    .Z(_1749_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5083_ (.A1(\mod.Data_Mem.F_M.MRAM[22][2] ),
    .A2(_1749_),
    .B(_1641_),
    .ZN(_1750_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5084_ (.I(_1524_),
    .Z(_1751_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5085_ (.I0(\mod.Data_Mem.F_M.MRAM[21][2] ),
    .I1(\mod.Data_Mem.F_M.MRAM[20][2] ),
    .S(_1701_),
    .Z(_1752_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5086_ (.A1(_1751_),
    .A2(_1752_),
    .ZN(_1753_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _5087_ (.A1(_1744_),
    .A2(_1748_),
    .B1(_1750_),
    .B2(_1753_),
    .C(_1616_),
    .ZN(_1754_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5088_ (.A1(_1508_),
    .A2(_1741_),
    .B(_1754_),
    .ZN(_1755_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5089_ (.I(_1499_),
    .Z(_1756_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5090_ (.I(_1756_),
    .Z(_1757_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5091_ (.A1(_1757_),
    .A2(\mod.Data_Mem.F_M.MRAM[31][2] ),
    .B1(_1721_),
    .B2(\mod.Data_Mem.F_M.MRAM[15][2] ),
    .ZN(_1758_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5092_ (.I(_1597_),
    .Z(_1759_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5093_ (.I0(_1755_),
    .I1(_1758_),
    .S(_1759_),
    .Z(_1760_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5094_ (.I0(\mod.Data_Mem.F_M.MRAM[775][2] ),
    .I1(\mod.Data_Mem.F_M.MRAM[774][2] ),
    .S(_1746_),
    .Z(_1761_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5095_ (.I0(\mod.Data_Mem.F_M.MRAM[773][2] ),
    .I1(\mod.Data_Mem.F_M.MRAM[772][2] ),
    .S(_1746_),
    .Z(_1762_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5096_ (.I0(_1761_),
    .I1(_1762_),
    .S(_1565_),
    .Z(_1763_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5097_ (.I(_1607_),
    .Z(_1764_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5098_ (.I(\mod.Data_Mem.F_M.MRAM[770][2] ),
    .ZN(_1765_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5099_ (.A1(_1708_),
    .A2(_1765_),
    .ZN(_1766_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5100_ (.A1(_1707_),
    .A2(\mod.Data_Mem.F_M.MRAM[771][2] ),
    .B(_1766_),
    .ZN(_1767_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5101_ (.A1(_1764_),
    .A2(_1767_),
    .ZN(_1768_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _5102_ (.I(_1701_),
    .Z(_1769_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5103_ (.I(\mod.Data_Mem.F_M.MRAM[768][2] ),
    .ZN(_1770_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5104_ (.A1(_1708_),
    .A2(_1770_),
    .ZN(_1771_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5105_ (.A1(_1769_),
    .A2(\mod.Data_Mem.F_M.MRAM[769][2] ),
    .B(_1771_),
    .ZN(_1772_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5106_ (.A1(_1603_),
    .A2(_1772_),
    .B(_1651_),
    .ZN(_1773_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5107_ (.A1(_1563_),
    .A2(_1763_),
    .B1(_1768_),
    .B2(_1773_),
    .ZN(_1774_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5108_ (.I(_1598_),
    .Z(_1775_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5109_ (.A1(\mod.Data_Mem.F_M.MRAM[783][2] ),
    .A2(_1775_),
    .ZN(_1776_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _5110_ (.A1(_1759_),
    .A2(_1774_),
    .B(_1776_),
    .C(_1508_),
    .ZN(_1777_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5111_ (.I(_1690_),
    .Z(_1778_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5112_ (.I(_1579_),
    .Z(_1779_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _5113_ (.A1(_1779_),
    .A2(\mod.Data_Mem.F_M.MRAM[790][2] ),
    .Z(_1780_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5114_ (.A1(_1778_),
    .A2(\mod.Data_Mem.F_M.MRAM[791][2] ),
    .B(_1780_),
    .ZN(_1781_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5115_ (.I(_1518_),
    .Z(_1782_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _5116_ (.I(_1567_),
    .Z(_1783_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5117_ (.I(\mod.Data_Mem.F_M.MRAM[788][2] ),
    .ZN(_1784_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5118_ (.A1(_1783_),
    .A2(_1784_),
    .ZN(_1785_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5119_ (.A1(_1782_),
    .A2(\mod.Data_Mem.F_M.MRAM[789][2] ),
    .B(_1785_),
    .ZN(_1786_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5120_ (.I(\mod.Data_Mem.F_M.MRAM[786][2] ),
    .ZN(_1787_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5121_ (.A1(_1715_),
    .A2(_1787_),
    .ZN(_1788_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5122_ (.A1(_1714_),
    .A2(\mod.Data_Mem.F_M.MRAM[787][2] ),
    .B(_1788_),
    .ZN(_1789_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5123_ (.I(_1513_),
    .Z(_1790_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5124_ (.I(_1790_),
    .Z(_1791_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5125_ (.I(\mod.Data_Mem.F_M.MRAM[784][2] ),
    .ZN(_1792_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5126_ (.A1(_1715_),
    .A2(_1792_),
    .ZN(_1793_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5127_ (.A1(_1791_),
    .A2(\mod.Data_Mem.F_M.MRAM[785][2] ),
    .B(_1793_),
    .ZN(_1794_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5128_ (.I(_1530_),
    .Z(_1795_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _5129_ (.I0(_1781_),
    .I1(_1786_),
    .I2(_1789_),
    .I3(_1794_),
    .S0(_1527_),
    .S1(_1795_),
    .Z(_1796_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5130_ (.A1(\mod.Data_Mem.F_M.MRAM[799][2] ),
    .A2(_1775_),
    .ZN(_1797_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _5131_ (.A1(_1759_),
    .A2(_1796_),
    .B(_1797_),
    .C(_1558_),
    .ZN(_1798_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5132_ (.I(_1669_),
    .Z(_1799_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _5133_ (.I(_1799_),
    .Z(_1800_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5134_ (.A1(_1777_),
    .A2(_1798_),
    .B(_1800_),
    .ZN(_1801_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _5135_ (.A1(_1729_),
    .A2(_1627_),
    .B1(_1760_),
    .B2(_1670_),
    .C(_1801_),
    .ZN(_0002_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5136_ (.I(_1695_),
    .Z(_1802_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5137_ (.A1(_1669_),
    .A2(_1626_),
    .ZN(_1803_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5138_ (.I(_1799_),
    .Z(_1804_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5139_ (.I(_1641_),
    .Z(_1805_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5140_ (.I0(\mod.Data_Mem.F_M.MRAM[21][3] ),
    .I1(\mod.Data_Mem.F_M.MRAM[20][3] ),
    .S(_1510_),
    .Z(_1806_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _5141_ (.A1(\mod.Data_Mem.F_M.MRAM[22][3] ),
    .A2(_1601_),
    .B1(_1730_),
    .B2(_1806_),
    .C(_1507_),
    .ZN(_1807_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5142_ (.I0(\mod.Data_Mem.F_M.MRAM[5][3] ),
    .I1(\mod.Data_Mem.F_M.MRAM[4][3] ),
    .S(_1510_),
    .Z(_1808_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5143_ (.I(_1543_),
    .Z(_1809_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _5144_ (.A1(\mod.Data_Mem.F_M.MRAM[6][3] ),
    .A2(_1645_),
    .B1(_1808_),
    .B2(_1809_),
    .C(_1557_),
    .ZN(_1810_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5145_ (.I(_1503_),
    .Z(_1811_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5146_ (.I(_1811_),
    .Z(_1812_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5147_ (.I(_1517_),
    .Z(_1813_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _5148_ (.I(_1813_),
    .Z(_1814_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _5149_ (.I0(\mod.Data_Mem.F_M.MRAM[3][3] ),
    .I1(\mod.Data_Mem.F_M.MRAM[1][3] ),
    .I2(\mod.Data_Mem.F_M.MRAM[0][3] ),
    .I3(\mod.Data_Mem.F_M.MRAM[2][3] ),
    .S0(_1812_),
    .S1(_1814_),
    .Z(_1815_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _5150_ (.I(_1586_),
    .Z(_1816_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5151_ (.I0(\mod.Data_Mem.F_M.MRAM[19][3] ),
    .I1(\mod.Data_Mem.F_M.MRAM[18][3] ),
    .S(_1816_),
    .Z(_1817_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5152_ (.A1(_1574_),
    .A2(_1817_),
    .ZN(_1818_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5153_ (.I0(\mod.Data_Mem.F_M.MRAM[17][3] ),
    .I1(\mod.Data_Mem.F_M.MRAM[16][3] ),
    .S(_1816_),
    .Z(_1819_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5154_ (.A1(_1584_),
    .A2(_1819_),
    .ZN(_1820_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _5155_ (.A1(_1557_),
    .A2(_1818_),
    .A3(_1820_),
    .ZN(_1821_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5156_ (.I(_1530_),
    .Z(_1822_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _5157_ (.A1(_1653_),
    .A2(_1815_),
    .B(_1821_),
    .C(_1822_),
    .ZN(_1823_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _5158_ (.A1(_1805_),
    .A2(_1807_),
    .A3(_1810_),
    .B(_1823_),
    .ZN(_1824_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5159_ (.A1(_1804_),
    .A2(_1824_),
    .ZN(_1825_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5160_ (.I(_1663_),
    .Z(_1826_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5161_ (.I0(\mod.Data_Mem.F_M.MRAM[785][3] ),
    .I1(\mod.Data_Mem.F_M.MRAM[784][3] ),
    .S(_1685_),
    .Z(_1827_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5162_ (.A1(_1826_),
    .A2(_1827_),
    .ZN(_1828_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _5163_ (.I(_1816_),
    .Z(_1829_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5164_ (.I0(\mod.Data_Mem.F_M.MRAM[787][3] ),
    .I1(\mod.Data_Mem.F_M.MRAM[786][3] ),
    .S(_1829_),
    .Z(_1830_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5165_ (.A1(_1608_),
    .A2(_1830_),
    .B(_1614_),
    .ZN(_1831_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5166_ (.I0(\mod.Data_Mem.F_M.MRAM[791][3] ),
    .I1(\mod.Data_Mem.F_M.MRAM[790][3] ),
    .S(_1581_),
    .Z(_1832_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5167_ (.A1(_1764_),
    .A2(_1832_),
    .B(_1531_),
    .ZN(_1833_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5168_ (.I(_1663_),
    .Z(_1834_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5169_ (.I(_1586_),
    .Z(_1835_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _5170_ (.I(_1835_),
    .Z(_1836_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5171_ (.I0(\mod.Data_Mem.F_M.MRAM[789][3] ),
    .I1(\mod.Data_Mem.F_M.MRAM[788][3] ),
    .S(_1836_),
    .Z(_1837_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5172_ (.A1(_1834_),
    .A2(_1837_),
    .ZN(_1838_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5173_ (.A1(_1828_),
    .A2(_1831_),
    .B1(_1833_),
    .B2(_1838_),
    .ZN(_1839_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5174_ (.I(_1690_),
    .Z(_1840_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _5175_ (.A1(_1835_),
    .A2(\mod.Data_Mem.F_M.MRAM[774][3] ),
    .Z(_1841_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5176_ (.A1(_1840_),
    .A2(\mod.Data_Mem.F_M.MRAM[775][3] ),
    .B(_1841_),
    .ZN(_1842_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5177_ (.A1(_1745_),
    .A2(_1842_),
    .ZN(_1843_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _5178_ (.I(_1526_),
    .Z(_1844_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5179_ (.I(_1578_),
    .Z(_1845_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5180_ (.I(\mod.Data_Mem.F_M.MRAM[772][3] ),
    .ZN(_1846_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5181_ (.A1(_1647_),
    .A2(_1846_),
    .ZN(_1847_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5182_ (.A1(_1845_),
    .A2(\mod.Data_Mem.F_M.MRAM[773][3] ),
    .B(_1847_),
    .ZN(_1848_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5183_ (.A1(_1844_),
    .A2(_1848_),
    .ZN(_1849_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _5184_ (.A1(_1614_),
    .A2(_1843_),
    .A3(_1849_),
    .ZN(_1850_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5185_ (.I(\mod.Data_Mem.F_M.MRAM[770][3] ),
    .ZN(_1851_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5186_ (.A1(_1647_),
    .A2(_1851_),
    .ZN(_1852_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5187_ (.A1(_1845_),
    .A2(\mod.Data_Mem.F_M.MRAM[771][3] ),
    .B(_1852_),
    .ZN(_1853_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5188_ (.A1(_1745_),
    .A2(_1853_),
    .ZN(_1854_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5189_ (.I(\mod.Data_Mem.F_M.MRAM[768][3] ),
    .ZN(_1855_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5190_ (.A1(_1658_),
    .A2(_1855_),
    .ZN(_1856_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5191_ (.A1(_1836_),
    .A2(\mod.Data_Mem.F_M.MRAM[769][3] ),
    .B(_1856_),
    .ZN(_1857_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5192_ (.A1(_1844_),
    .A2(_1857_),
    .ZN(_1858_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _5193_ (.A1(_1642_),
    .A2(_1854_),
    .A3(_1858_),
    .ZN(_1859_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _5194_ (.A1(_1721_),
    .A2(_1850_),
    .A3(_1859_),
    .ZN(_1860_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _5195_ (.A1(_1621_),
    .A2(_1839_),
    .B(_1860_),
    .C(_1490_),
    .ZN(_1861_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _5196_ (.A1(_1552_),
    .A2(_1825_),
    .A3(_1861_),
    .ZN(_1862_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5197_ (.I(_1557_),
    .Z(_1863_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5198_ (.A1(\mod.Data_Mem.F_M.MRAM[783][3] ),
    .A2(_1863_),
    .ZN(_1864_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5199_ (.A1(\mod.Data_Mem.F_M.MRAM[799][3] ),
    .A2(_1621_),
    .B(_1625_),
    .ZN(_1865_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5200_ (.I(_1669_),
    .Z(_1866_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _5201_ (.A1(_1757_),
    .A2(\mod.Data_Mem.F_M.MRAM[15][3] ),
    .B1(\mod.Data_Mem.F_M.MRAM[31][3] ),
    .B2(_1721_),
    .C(_1866_),
    .ZN(_1867_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _5202_ (.A1(_1864_),
    .A2(_1865_),
    .B(_1867_),
    .C(_1699_),
    .ZN(_1868_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _5203_ (.A1(_1631_),
    .A2(_1862_),
    .A3(_1868_),
    .ZN(_1869_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5204_ (.A1(_1802_),
    .A2(_1803_),
    .B(_1869_),
    .ZN(_0003_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5205_ (.I(\mod.Data_Mem.F_M.MRAM[15][4] ),
    .Z(_1870_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5206_ (.A1(_1870_),
    .A2(_1673_),
    .ZN(_1871_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5207_ (.I(_1550_),
    .Z(_1872_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _5208_ (.I(_1587_),
    .Z(_1873_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5209_ (.I0(\mod.Data_Mem.F_M.MRAM[5][4] ),
    .I1(\mod.Data_Mem.F_M.MRAM[4][4] ),
    .S(_1873_),
    .Z(_1874_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5210_ (.I(_1646_),
    .Z(_1875_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5211_ (.I0(\mod.Data_Mem.F_M.MRAM[7][4] ),
    .I1(\mod.Data_Mem.F_M.MRAM[6][4] ),
    .S(_1875_),
    .Z(_1876_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _5212_ (.I(_1580_),
    .Z(_1877_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5213_ (.I0(\mod.Data_Mem.F_M.MRAM[1][4] ),
    .I1(\mod.Data_Mem.F_M.MRAM[0][4] ),
    .S(_1877_),
    .Z(_1878_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5214_ (.I(_1790_),
    .Z(_1879_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5215_ (.I0(\mod.Data_Mem.F_M.MRAM[3][4] ),
    .I1(\mod.Data_Mem.F_M.MRAM[2][4] ),
    .S(_1879_),
    .Z(_1880_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _5216_ (.I(_1607_),
    .Z(_1881_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5217_ (.I(_1530_),
    .Z(_1882_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _5218_ (.I0(_1874_),
    .I1(_1876_),
    .I2(_1878_),
    .I3(_1880_),
    .S0(_1881_),
    .S1(_1882_),
    .Z(_1883_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5219_ (.I(_1653_),
    .Z(_1884_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5220_ (.A1(_1872_),
    .A2(_1883_),
    .B(_1884_),
    .ZN(_1885_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5221_ (.I(_1672_),
    .Z(_1886_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5222_ (.A1(\mod.Data_Mem.F_M.MRAM[31][4] ),
    .A2(_1886_),
    .ZN(_1887_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5223_ (.I(_1550_),
    .Z(_1888_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5224_ (.I0(\mod.Data_Mem.F_M.MRAM[23][4] ),
    .I1(\mod.Data_Mem.F_M.MRAM[22][4] ),
    .S(_1588_),
    .Z(_1889_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _5225_ (.I(_1587_),
    .Z(_1890_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5226_ (.I0(\mod.Data_Mem.F_M.MRAM[21][4] ),
    .I1(\mod.Data_Mem.F_M.MRAM[20][4] ),
    .S(_1890_),
    .Z(_1891_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _5227_ (.I(_1790_),
    .Z(_1892_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5228_ (.I0(\mod.Data_Mem.F_M.MRAM[19][4] ),
    .I1(\mod.Data_Mem.F_M.MRAM[18][4] ),
    .S(_1892_),
    .Z(_1893_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _5229_ (.I(_1813_),
    .Z(_1894_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5230_ (.I0(\mod.Data_Mem.F_M.MRAM[17][4] ),
    .I1(\mod.Data_Mem.F_M.MRAM[16][4] ),
    .S(_1894_),
    .Z(_1895_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _5231_ (.I0(_1889_),
    .I1(_1891_),
    .I2(_1893_),
    .I3(_1895_),
    .S0(_1751_),
    .S1(_1882_),
    .Z(_1896_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5232_ (.A1(_1888_),
    .A2(_1896_),
    .B(_1633_),
    .ZN(_1897_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5233_ (.I(_1799_),
    .Z(_1898_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5234_ (.A1(_1898_),
    .A2(_1628_),
    .ZN(_1899_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _5235_ (.A1(_1871_),
    .A2(_1885_),
    .B1(_1887_),
    .B2(_1897_),
    .C(_1899_),
    .ZN(_1900_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5236_ (.I(\mod.Data_Mem.F_M.MRAM[783][4] ),
    .Z(_1901_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5237_ (.A1(_1901_),
    .A2(_1699_),
    .ZN(_1902_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5238_ (.I(_1813_),
    .Z(_1903_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5239_ (.I0(\mod.Data_Mem.F_M.MRAM[773][4] ),
    .I1(\mod.Data_Mem.F_M.MRAM[772][4] ),
    .S(_1903_),
    .Z(_1904_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5240_ (.I0(\mod.Data_Mem.F_M.MRAM[775][4] ),
    .I1(\mod.Data_Mem.F_M.MRAM[774][4] ),
    .S(_1836_),
    .Z(_1905_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _5241_ (.I(_1835_),
    .Z(_1906_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5242_ (.I0(\mod.Data_Mem.F_M.MRAM[769][4] ),
    .I1(\mod.Data_Mem.F_M.MRAM[768][4] ),
    .S(_1906_),
    .Z(_1907_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _5243_ (.I(_1587_),
    .Z(_1908_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5244_ (.I0(\mod.Data_Mem.F_M.MRAM[771][4] ),
    .I1(\mod.Data_Mem.F_M.MRAM[770][4] ),
    .S(_1908_),
    .Z(_1909_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _5245_ (.I(_1644_),
    .Z(_1910_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _5246_ (.I0(_1904_),
    .I1(_1905_),
    .I2(_1907_),
    .I3(_1909_),
    .S0(_1910_),
    .S1(_1805_),
    .Z(_1911_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5247_ (.A1(_1552_),
    .A2(_1911_),
    .B(_1884_),
    .ZN(_1912_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5248_ (.I(_1672_),
    .Z(_1913_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5249_ (.I(_1503_),
    .Z(_1914_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5250_ (.I(_1914_),
    .Z(_1915_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _5251_ (.I0(\mod.Data_Mem.F_M.MRAM[791][4] ),
    .I1(\mod.Data_Mem.F_M.MRAM[788][4] ),
    .I2(\mod.Data_Mem.F_M.MRAM[789][4] ),
    .I3(\mod.Data_Mem.F_M.MRAM[790][4] ),
    .S0(_1829_),
    .S1(_1915_),
    .Z(_1916_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5252_ (.A1(_1700_),
    .A2(_1916_),
    .ZN(_1917_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _5253_ (.I(_1779_),
    .Z(_1918_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5254_ (.I(\mod.Data_Mem.F_M.MRAM[787][4] ),
    .ZN(_1919_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5255_ (.A1(_1906_),
    .A2(\mod.Data_Mem.F_M.MRAM[786][4] ),
    .ZN(_1920_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5256_ (.A1(_1918_),
    .A2(_1919_),
    .B(_1920_),
    .ZN(_1921_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5257_ (.I0(\mod.Data_Mem.F_M.MRAM[785][4] ),
    .I1(\mod.Data_Mem.F_M.MRAM[784][4] ),
    .S(_1580_),
    .Z(_1922_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _5258_ (.A1(_1704_),
    .A2(_1922_),
    .Z(_1923_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _5259_ (.A1(_1834_),
    .A2(_1921_),
    .B(_1923_),
    .C(_1642_),
    .ZN(_1924_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5260_ (.A1(_1917_),
    .A2(_1924_),
    .B(_1674_),
    .ZN(_1925_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5261_ (.A1(\mod.Data_Mem.F_M.MRAM[799][4] ),
    .A2(_1913_),
    .B(_1925_),
    .ZN(_1926_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5262_ (.I(_1653_),
    .Z(_1927_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _5263_ (.A1(_1902_),
    .A2(_1912_),
    .B1(_1926_),
    .B2(_1927_),
    .C(_1629_),
    .ZN(_1928_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _5264_ (.A1(_1900_),
    .A2(_1928_),
    .Z(_1929_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5265_ (.I(_1929_),
    .Z(_0004_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5266_ (.A1(\mod.Data_Mem.F_M.MRAM[799][5] ),
    .A2(_1599_),
    .ZN(_1930_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5267_ (.I(_1695_),
    .Z(_1931_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5268_ (.I(_1890_),
    .Z(_1932_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5269_ (.I(_1692_),
    .Z(_1933_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5270_ (.I(\mod.Data_Mem.F_M.MRAM[788][5] ),
    .ZN(_1934_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5271_ (.A1(_1933_),
    .A2(_1934_),
    .ZN(_1935_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5272_ (.A1(_1932_),
    .A2(\mod.Data_Mem.F_M.MRAM[789][5] ),
    .B(_1935_),
    .ZN(_1936_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5273_ (.I0(\mod.Data_Mem.F_M.MRAM[791][5] ),
    .I1(\mod.Data_Mem.F_M.MRAM[790][5] ),
    .S(_1783_),
    .Z(_1937_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5274_ (.A1(_1645_),
    .A2(_1937_),
    .ZN(_1938_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _5275_ (.A1(_1931_),
    .A2(_1936_),
    .B(_1938_),
    .C(_1563_),
    .ZN(_1939_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5276_ (.I(_1573_),
    .Z(_1940_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5277_ (.I(_1940_),
    .Z(_1941_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _5278_ (.I(_1514_),
    .Z(_1942_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5279_ (.I0(\mod.Data_Mem.F_M.MRAM[787][5] ),
    .I1(\mod.Data_Mem.F_M.MRAM[786][5] ),
    .S(_1942_),
    .Z(_1943_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5280_ (.A1(_1941_),
    .A2(_1943_),
    .ZN(_1944_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5281_ (.I0(\mod.Data_Mem.F_M.MRAM[785][5] ),
    .I1(\mod.Data_Mem.F_M.MRAM[784][5] ),
    .S(_1942_),
    .Z(_1945_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5282_ (.A1(_1826_),
    .A2(_1945_),
    .ZN(_1946_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _5283_ (.A1(_1805_),
    .A2(_1944_),
    .A3(_1946_),
    .ZN(_1947_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _5284_ (.A1(_1551_),
    .A2(_1939_),
    .A3(_1947_),
    .ZN(_1948_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _5285_ (.A1(_1927_),
    .A2(_1930_),
    .A3(_1948_),
    .ZN(_1949_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5286_ (.I0(\mod.Data_Mem.F_M.MRAM[773][5] ),
    .I1(\mod.Data_Mem.F_M.MRAM[772][5] ),
    .S(_1612_),
    .Z(_1950_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5287_ (.I(_1816_),
    .Z(_1951_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5288_ (.I0(\mod.Data_Mem.F_M.MRAM[775][5] ),
    .I1(\mod.Data_Mem.F_M.MRAM[774][5] ),
    .S(_1951_),
    .Z(_1952_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5289_ (.I(_1579_),
    .Z(_1953_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _5290_ (.I(_1953_),
    .Z(_1954_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5291_ (.I(\mod.Data_Mem.F_M.MRAM[769][5] ),
    .ZN(_1955_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5292_ (.A1(_1875_),
    .A2(\mod.Data_Mem.F_M.MRAM[768][5] ),
    .ZN(_1956_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5293_ (.A1(_1954_),
    .A2(_1955_),
    .B(_1956_),
    .ZN(_1957_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5294_ (.I0(\mod.Data_Mem.F_M.MRAM[771][5] ),
    .I1(\mod.Data_Mem.F_M.MRAM[770][5] ),
    .S(_1783_),
    .Z(_1958_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _5295_ (.I0(_1950_),
    .I1(_1952_),
    .I2(_1957_),
    .I3(_1958_),
    .S0(_1745_),
    .S1(_1822_),
    .Z(_1959_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5296_ (.A1(_1622_),
    .A2(_1959_),
    .ZN(_1960_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5297_ (.A1(\mod.Data_Mem.F_M.MRAM[783][5] ),
    .A2(_1599_),
    .ZN(_1961_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _5298_ (.A1(_1633_),
    .A2(_1960_),
    .A3(_1961_),
    .ZN(_1962_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _5299_ (.A1(_1631_),
    .A2(_1949_),
    .A3(_1962_),
    .ZN(_1963_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _5300_ (.I(_1724_),
    .Z(_1964_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5301_ (.I(_1964_),
    .Z(_1965_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5302_ (.I(_1965_),
    .Z(_1966_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5303_ (.A1(\mod.Data_Mem.F_M.MRAM[15][5] ),
    .A2(_1599_),
    .ZN(_1967_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _5304_ (.I(_1509_),
    .Z(_1968_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5305_ (.I0(\mod.Data_Mem.F_M.MRAM[5][5] ),
    .I1(\mod.Data_Mem.F_M.MRAM[4][5] ),
    .S(_1968_),
    .Z(_1969_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5306_ (.I0(\mod.Data_Mem.F_M.MRAM[7][5] ),
    .I1(\mod.Data_Mem.F_M.MRAM[6][5] ),
    .S(_1515_),
    .Z(_1970_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5307_ (.I(\mod.Data_Mem.F_M.MRAM[1][5] ),
    .ZN(_1971_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5308_ (.A1(_1942_),
    .A2(\mod.Data_Mem.F_M.MRAM[0][5] ),
    .ZN(_1972_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5309_ (.A1(_1769_),
    .A2(_1971_),
    .B(_1972_),
    .ZN(_1973_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5310_ (.I0(\mod.Data_Mem.F_M.MRAM[3][5] ),
    .I1(\mod.Data_Mem.F_M.MRAM[2][5] ),
    .S(_1968_),
    .Z(_1974_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _5311_ (.I0(_1969_),
    .I1(_1970_),
    .I2(_1973_),
    .I3(_1974_),
    .S0(_1695_),
    .S1(_1795_),
    .Z(_1975_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5312_ (.A1(_1622_),
    .A2(_1975_),
    .B(_1863_),
    .ZN(_1976_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5313_ (.A1(\mod.Data_Mem.F_M.MRAM[31][5] ),
    .A2(_1759_),
    .ZN(_1977_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5314_ (.I0(\mod.Data_Mem.F_M.MRAM[23][5] ),
    .I1(\mod.Data_Mem.F_M.MRAM[22][5] ),
    .S(_1568_),
    .Z(_1978_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5315_ (.I0(\mod.Data_Mem.F_M.MRAM[21][5] ),
    .I1(\mod.Data_Mem.F_M.MRAM[20][5] ),
    .S(_1968_),
    .Z(_1979_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5316_ (.I0(\mod.Data_Mem.F_M.MRAM[19][5] ),
    .I1(\mod.Data_Mem.F_M.MRAM[18][5] ),
    .S(_1681_),
    .Z(_1980_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5317_ (.I0(\mod.Data_Mem.F_M.MRAM[17][5] ),
    .I1(\mod.Data_Mem.F_M.MRAM[16][5] ),
    .S(_1568_),
    .Z(_1981_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _5318_ (.I0(_1978_),
    .I1(_1979_),
    .I2(_1980_),
    .I3(_1981_),
    .S0(_1527_),
    .S1(_1795_),
    .Z(_1982_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5319_ (.A1(_1551_),
    .A2(_1982_),
    .B(_1508_),
    .ZN(_1983_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5320_ (.A1(_1967_),
    .A2(_1976_),
    .B1(_1977_),
    .B2(_1983_),
    .ZN(_1984_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5321_ (.A1(_1966_),
    .A2(_1984_),
    .ZN(_1985_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5322_ (.A1(_1899_),
    .A2(_1963_),
    .B(_1985_),
    .ZN(_0005_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5323_ (.A1(\mod.Data_Mem.F_M.MRAM[15][6] ),
    .A2(_1673_),
    .ZN(_1986_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5324_ (.I0(\mod.Data_Mem.F_M.MRAM[5][6] ),
    .I1(\mod.Data_Mem.F_M.MRAM[4][6] ),
    .S(_1873_),
    .Z(_1987_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5325_ (.I0(\mod.Data_Mem.F_M.MRAM[7][6] ),
    .I1(\mod.Data_Mem.F_M.MRAM[6][6] ),
    .S(_1873_),
    .Z(_1988_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5326_ (.I0(\mod.Data_Mem.F_M.MRAM[1][6] ),
    .I1(\mod.Data_Mem.F_M.MRAM[0][6] ),
    .S(_1609_),
    .Z(_1989_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5327_ (.I0(\mod.Data_Mem.F_M.MRAM[3][6] ),
    .I1(\mod.Data_Mem.F_M.MRAM[2][6] ),
    .S(_1877_),
    .Z(_1990_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _5328_ (.I0(_1987_),
    .I1(_1988_),
    .I2(_1989_),
    .I3(_1990_),
    .S0(_1881_),
    .S1(_1882_),
    .Z(_1991_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5329_ (.A1(_1872_),
    .A2(_1991_),
    .B(_1863_),
    .ZN(_1992_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5330_ (.A1(\mod.Data_Mem.F_M.MRAM[31][6] ),
    .A2(_1886_),
    .ZN(_1993_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5331_ (.I0(\mod.Data_Mem.F_M.MRAM[23][6] ),
    .I1(\mod.Data_Mem.F_M.MRAM[22][6] ),
    .S(_1708_),
    .Z(_1994_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5332_ (.I0(\mod.Data_Mem.F_M.MRAM[21][6] ),
    .I1(\mod.Data_Mem.F_M.MRAM[20][6] ),
    .S(_1892_),
    .Z(_1995_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5333_ (.I0(\mod.Data_Mem.F_M.MRAM[19][6] ),
    .I1(\mod.Data_Mem.F_M.MRAM[18][6] ),
    .S(_1892_),
    .Z(_1996_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5334_ (.I0(\mod.Data_Mem.F_M.MRAM[17][6] ),
    .I1(\mod.Data_Mem.F_M.MRAM[16][6] ),
    .S(_1894_),
    .Z(_1997_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _5335_ (.I0(_1994_),
    .I1(_1995_),
    .I2(_1996_),
    .I3(_1997_),
    .S0(_1844_),
    .S1(_1882_),
    .Z(_1998_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5336_ (.A1(_1888_),
    .A2(_1998_),
    .B(_1633_),
    .ZN(_1999_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _5337_ (.A1(_1986_),
    .A2(_1992_),
    .B1(_1993_),
    .B2(_1999_),
    .C(_1899_),
    .ZN(_2000_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5338_ (.A1(\mod.Data_Mem.F_M.MRAM[783][6] ),
    .A2(_1699_),
    .ZN(_2001_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5339_ (.I0(\mod.Data_Mem.F_M.MRAM[769][6] ),
    .I1(\mod.Data_Mem.F_M.MRAM[768][6] ),
    .S(_1814_),
    .Z(_2002_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5340_ (.I0(\mod.Data_Mem.F_M.MRAM[771][6] ),
    .I1(\mod.Data_Mem.F_M.MRAM[770][6] ),
    .S(_1836_),
    .Z(_2003_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5341_ (.I0(\mod.Data_Mem.F_M.MRAM[773][6] ),
    .I1(\mod.Data_Mem.F_M.MRAM[772][6] ),
    .S(_1906_),
    .Z(_2004_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5342_ (.I0(\mod.Data_Mem.F_M.MRAM[775][6] ),
    .I1(\mod.Data_Mem.F_M.MRAM[774][6] ),
    .S(_1908_),
    .Z(_2005_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _5343_ (.I0(_2002_),
    .I1(_2003_),
    .I2(_2004_),
    .I3(_2005_),
    .S0(_1910_),
    .S1(_1590_),
    .Z(_2006_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5344_ (.A1(_1872_),
    .A2(_2006_),
    .B(_1884_),
    .ZN(_2007_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5345_ (.I(_1914_),
    .Z(_2008_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5346_ (.I(_2008_),
    .Z(_2009_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _5347_ (.I0(\mod.Data_Mem.F_M.MRAM[791][6] ),
    .I1(\mod.Data_Mem.F_M.MRAM[788][6] ),
    .I2(\mod.Data_Mem.F_M.MRAM[789][6] ),
    .I3(\mod.Data_Mem.F_M.MRAM[790][6] ),
    .S0(_1829_),
    .S1(_2009_),
    .Z(_2010_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5348_ (.A1(_1700_),
    .A2(_2010_),
    .ZN(_2011_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5349_ (.I(_1602_),
    .Z(_2012_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5350_ (.I(\mod.Data_Mem.F_M.MRAM[787][6] ),
    .ZN(_2013_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5351_ (.A1(_1903_),
    .A2(\mod.Data_Mem.F_M.MRAM[786][6] ),
    .ZN(_2014_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5352_ (.A1(_1933_),
    .A2(_2013_),
    .B(_2014_),
    .ZN(_2015_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5353_ (.I0(\mod.Data_Mem.F_M.MRAM[785][6] ),
    .I1(\mod.Data_Mem.F_M.MRAM[784][6] ),
    .S(_1580_),
    .Z(_2016_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _5354_ (.A1(_1704_),
    .A2(_2016_),
    .Z(_2017_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _5355_ (.A1(_2012_),
    .A2(_2015_),
    .B(_2017_),
    .C(_1822_),
    .ZN(_2018_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5356_ (.A1(_2011_),
    .A2(_2018_),
    .B(_1775_),
    .ZN(_2019_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5357_ (.A1(\mod.Data_Mem.F_M.MRAM[799][6] ),
    .A2(_1913_),
    .B(_2019_),
    .ZN(_2020_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _5358_ (.A1(_2001_),
    .A2(_2007_),
    .B1(_2020_),
    .B2(_1927_),
    .C(_1629_),
    .ZN(_2021_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _5359_ (.A1(_2000_),
    .A2(_2021_),
    .Z(_2022_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5360_ (.I(_2022_),
    .Z(_0006_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5361_ (.A1(\mod.Data_Mem.F_M.MRAM[15][7] ),
    .A2(_1886_),
    .ZN(_2023_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5362_ (.I0(\mod.Data_Mem.F_M.MRAM[1][7] ),
    .I1(\mod.Data_Mem.F_M.MRAM[0][7] ),
    .S(_1879_),
    .Z(_2024_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _5363_ (.I(_1835_),
    .Z(_2025_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5364_ (.I0(\mod.Data_Mem.F_M.MRAM[3][7] ),
    .I1(\mod.Data_Mem.F_M.MRAM[2][7] ),
    .S(_2025_),
    .Z(_2026_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5365_ (.I0(\mod.Data_Mem.F_M.MRAM[5][7] ),
    .I1(\mod.Data_Mem.F_M.MRAM[4][7] ),
    .S(_1877_),
    .Z(_2027_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5366_ (.I0(\mod.Data_Mem.F_M.MRAM[7][7] ),
    .I1(\mod.Data_Mem.F_M.MRAM[6][7] ),
    .S(_1877_),
    .Z(_2028_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _5367_ (.I0(_2024_),
    .I1(_2026_),
    .I2(_2027_),
    .I3(_2028_),
    .S0(_1881_),
    .S1(_1590_),
    .Z(_2029_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5368_ (.A1(_1888_),
    .A2(_2029_),
    .B(_1863_),
    .ZN(_2030_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5369_ (.A1(\mod.Data_Mem.F_M.MRAM[31][7] ),
    .A2(_1913_),
    .ZN(_2031_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5370_ (.I0(\mod.Data_Mem.F_M.MRAM[23][7] ),
    .I1(\mod.Data_Mem.F_M.MRAM[22][7] ),
    .S(_1588_),
    .Z(_2032_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5371_ (.I0(\mod.Data_Mem.F_M.MRAM[21][7] ),
    .I1(\mod.Data_Mem.F_M.MRAM[20][7] ),
    .S(_1890_),
    .Z(_2033_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5372_ (.I0(\mod.Data_Mem.F_M.MRAM[19][7] ),
    .I1(\mod.Data_Mem.F_M.MRAM[18][7] ),
    .S(_1892_),
    .Z(_2034_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5373_ (.I0(\mod.Data_Mem.F_M.MRAM[17][7] ),
    .I1(\mod.Data_Mem.F_M.MRAM[16][7] ),
    .S(_1894_),
    .Z(_2035_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _5374_ (.I0(_2032_),
    .I1(_2033_),
    .I2(_2034_),
    .I3(_2035_),
    .S0(_1844_),
    .S1(_1642_),
    .Z(_2036_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5375_ (.A1(_1888_),
    .A2(_2036_),
    .B(_1621_),
    .ZN(_2037_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _5376_ (.A1(_2023_),
    .A2(_2030_),
    .B1(_2031_),
    .B2(_2037_),
    .C(_1899_),
    .ZN(_2038_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5377_ (.A1(\mod.Data_Mem.F_M.MRAM[783][7] ),
    .A2(_1673_),
    .ZN(_2039_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5378_ (.I0(\mod.Data_Mem.F_M.MRAM[769][7] ),
    .I1(\mod.Data_Mem.F_M.MRAM[768][7] ),
    .S(_1814_),
    .Z(_2040_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5379_ (.I0(\mod.Data_Mem.F_M.MRAM[771][7] ),
    .I1(\mod.Data_Mem.F_M.MRAM[770][7] ),
    .S(_1903_),
    .Z(_2041_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5380_ (.I0(\mod.Data_Mem.F_M.MRAM[773][7] ),
    .I1(\mod.Data_Mem.F_M.MRAM[772][7] ),
    .S(_1906_),
    .Z(_2042_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5381_ (.I0(\mod.Data_Mem.F_M.MRAM[775][7] ),
    .I1(\mod.Data_Mem.F_M.MRAM[774][7] ),
    .S(_1908_),
    .Z(_2043_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _5382_ (.I(_1607_),
    .Z(_2044_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _5383_ (.I0(_2040_),
    .I1(_2041_),
    .I2(_2042_),
    .I3(_2043_),
    .S0(_2044_),
    .S1(_1590_),
    .Z(_2045_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5384_ (.A1(_1872_),
    .A2(_2045_),
    .B(_1884_),
    .ZN(_2046_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _5385_ (.I0(\mod.Data_Mem.F_M.MRAM[791][7] ),
    .I1(\mod.Data_Mem.F_M.MRAM[788][7] ),
    .I2(\mod.Data_Mem.F_M.MRAM[789][7] ),
    .I3(\mod.Data_Mem.F_M.MRAM[790][7] ),
    .S0(_1829_),
    .S1(_2009_),
    .Z(_2047_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5386_ (.A1(_1700_),
    .A2(_2047_),
    .ZN(_2048_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5387_ (.I(\mod.Data_Mem.F_M.MRAM[787][7] ),
    .ZN(_2049_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5388_ (.A1(_1875_),
    .A2(\mod.Data_Mem.F_M.MRAM[786][7] ),
    .ZN(_2050_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5389_ (.A1(_1918_),
    .A2(_2049_),
    .B(_2050_),
    .ZN(_2051_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5390_ (.I0(\mod.Data_Mem.F_M.MRAM[785][7] ),
    .I1(\mod.Data_Mem.F_M.MRAM[784][7] ),
    .S(_1813_),
    .Z(_2052_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _5391_ (.A1(_1704_),
    .A2(_2052_),
    .Z(_2053_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _5392_ (.A1(_2012_),
    .A2(_2051_),
    .B(_2053_),
    .C(_1822_),
    .ZN(_2054_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5393_ (.A1(_2048_),
    .A2(_2054_),
    .B(_1775_),
    .ZN(_2055_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5394_ (.A1(\mod.Data_Mem.F_M.MRAM[799][7] ),
    .A2(_1913_),
    .B(_2055_),
    .ZN(_2056_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _5395_ (.A1(_2039_),
    .A2(_2046_),
    .B1(_2056_),
    .B2(_1927_),
    .C(_1629_),
    .ZN(_2057_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _5396_ (.A1(_2038_),
    .A2(_2057_),
    .Z(_2058_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5397_ (.I(_2058_),
    .Z(_0007_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5398_ (.I(_1522_),
    .Z(_2059_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5399_ (.I(_2059_),
    .Z(_2060_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5400_ (.I(_2060_),
    .Z(_2061_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5401_ (.I(_2061_),
    .Z(_2062_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5402_ (.I(_2062_),
    .Z(_2063_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5403_ (.I(_1501_),
    .Z(_2064_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5404_ (.A1(_2064_),
    .A2(_1553_),
    .ZN(_2065_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5405_ (.A1(_1724_),
    .A2(_2065_),
    .ZN(_2066_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5406_ (.I(_2066_),
    .Z(_2067_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5407_ (.I(_2067_),
    .Z(_2068_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5408_ (.I(_2068_),
    .Z(_0010_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5409_ (.A1(_2063_),
    .A2(_0010_),
    .ZN(_0008_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5410_ (.I(_1595_),
    .Z(_2069_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5411_ (.I(_2069_),
    .Z(_2070_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5412_ (.I(_2070_),
    .Z(_2071_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5413_ (.I(_2071_),
    .Z(_2072_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5414_ (.I(_1725_),
    .Z(_2073_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5415_ (.I(_2073_),
    .Z(_2074_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5416_ (.I(_2065_),
    .Z(_2075_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5417_ (.I(_2075_),
    .Z(_2076_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5418_ (.I(_2076_),
    .Z(_2077_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _5419_ (.A1(_2072_),
    .A2(_2074_),
    .A3(_2077_),
    .ZN(_0009_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5420_ (.I(_1489_),
    .Z(_2078_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5421_ (.I(_2078_),
    .Z(_2079_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5422_ (.I(_2079_),
    .Z(_2080_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5423_ (.A1(_2080_),
    .A2(_2077_),
    .ZN(_0011_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5424_ (.I(_1701_),
    .Z(_2081_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5425_ (.A1(_2081_),
    .A2(_0010_),
    .ZN(_0016_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5426_ (.I(_2067_),
    .Z(_2082_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _5427_ (.A1(_1802_),
    .A2(_2082_),
    .Z(_2083_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5428_ (.I(_2083_),
    .Z(_0017_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5429_ (.I(_1725_),
    .Z(_2084_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5430_ (.I(_2084_),
    .Z(_2085_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5431_ (.I(_1549_),
    .Z(_2086_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5432_ (.I(_2086_),
    .Z(_2087_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _5433_ (.A1(_2085_),
    .A2(_2087_),
    .A3(_2076_),
    .ZN(_0018_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5434_ (.A1(_2080_),
    .A2(_2077_),
    .ZN(_0019_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5435_ (.A1(_2063_),
    .A2(_0010_),
    .ZN(_0024_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5436_ (.I(_2069_),
    .Z(_2088_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5437_ (.I(_2088_),
    .Z(_2089_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5438_ (.A1(_2089_),
    .A2(_2067_),
    .ZN(_2090_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5439_ (.I(_2090_),
    .ZN(_0025_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _5440_ (.A1(_2072_),
    .A2(_2074_),
    .A3(_2076_),
    .ZN(_0026_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5441_ (.A1(_2080_),
    .A2(_2077_),
    .ZN(_0027_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5442_ (.I(_2008_),
    .Z(_2091_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5443_ (.I(_1548_),
    .Z(_2092_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _5444_ (.A1(_2092_),
    .A2(_1619_),
    .ZN(_2093_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5445_ (.A1(_2078_),
    .A2(_2093_),
    .ZN(_2094_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5446_ (.A1(_2091_),
    .A2(_2094_),
    .ZN(_2095_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5447_ (.I(_1522_),
    .Z(_2096_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5448_ (.I(_2096_),
    .Z(_2097_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _5449_ (.A1(_1951_),
    .A2(\mod.Data_Mem.F_M.MRAM[799][0] ),
    .Z(_2098_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _5450_ (.A1(_2097_),
    .A2(\mod.Data_Mem.F_M.MRAM[798][0] ),
    .B(_2098_),
    .ZN(_2099_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5451_ (.I(_1535_),
    .Z(_2100_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5452_ (.A1(_2008_),
    .A2(_1554_),
    .ZN(_2101_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5453_ (.I(_2101_),
    .Z(_2102_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5454_ (.I(_2102_),
    .Z(_2103_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5455_ (.A1(_2100_),
    .A2(_2103_),
    .ZN(_2104_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5456_ (.A1(_2081_),
    .A2(_2104_),
    .ZN(_2105_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5457_ (.I(_1495_),
    .Z(_2106_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5458_ (.I(_2106_),
    .Z(_2107_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5459_ (.I(_2107_),
    .Z(_2108_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5460_ (.A1(_2069_),
    .A2(_2064_),
    .ZN(_2109_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5461_ (.I(_2109_),
    .Z(_2110_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5462_ (.A1(_2108_),
    .A2(_2110_),
    .ZN(_2111_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5463_ (.I0(\mod.Data_Mem.F_M.MRAM[30][0] ),
    .I1(\mod.Data_Mem.F_M.MRAM[31][0] ),
    .S(_1873_),
    .Z(_2112_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5464_ (.I(_1803_),
    .ZN(_2113_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5465_ (.A1(_2113_),
    .A2(_2066_),
    .ZN(_2114_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5466_ (.A1(_2111_),
    .A2(_2112_),
    .B(_2114_),
    .ZN(_2115_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5467_ (.A1(_2095_),
    .A2(_2099_),
    .B1(_2105_),
    .B2(_2115_),
    .ZN(_0032_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5468_ (.I(_1812_),
    .Z(_2116_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5469_ (.A1(_2116_),
    .A2(_1626_),
    .ZN(_2117_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5470_ (.I(_2117_),
    .Z(_2118_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5471_ (.I(_2090_),
    .Z(_2119_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _5472_ (.A1(_1951_),
    .A2(\mod.Data_Mem.F_M.MRAM[31][1] ),
    .Z(_2120_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5473_ (.A1(_2097_),
    .A2(\mod.Data_Mem.F_M.MRAM[30][1] ),
    .B(_2120_),
    .ZN(_2121_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5474_ (.I0(\mod.Data_Mem.F_M.MRAM[798][1] ),
    .I1(\mod.Data_Mem.F_M.MRAM[799][1] ),
    .S(_1908_),
    .Z(_2122_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5475_ (.A1(_2095_),
    .A2(_2122_),
    .ZN(_2123_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _5476_ (.A1(_2074_),
    .A2(_2118_),
    .B1(_2119_),
    .B2(_2121_),
    .C(_2123_),
    .ZN(_0033_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5477_ (.I0(\mod.Data_Mem.F_M.MRAM[30][2] ),
    .I1(\mod.Data_Mem.F_M.MRAM[31][2] ),
    .S(_1510_),
    .Z(_2124_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5478_ (.I0(\mod.Data_Mem.F_M.MRAM[798][2] ),
    .I1(\mod.Data_Mem.F_M.MRAM[799][2] ),
    .S(_1890_),
    .Z(_2125_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5479_ (.A1(_0025_),
    .A2(_2124_),
    .B1(_2125_),
    .B2(_2095_),
    .ZN(_2126_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5480_ (.A1(_1803_),
    .A2(_2126_),
    .ZN(_0034_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5481_ (.I0(\mod.Data_Mem.F_M.MRAM[30][3] ),
    .I1(\mod.Data_Mem.F_M.MRAM[31][3] ),
    .S(_1845_),
    .Z(_2127_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5482_ (.A1(_2110_),
    .A2(_2127_),
    .ZN(_2128_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5483_ (.I(_2096_),
    .Z(_2129_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _5484_ (.A1(_1879_),
    .A2(\mod.Data_Mem.F_M.MRAM[798][3] ),
    .Z(_2130_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5485_ (.A1(_2129_),
    .A2(\mod.Data_Mem.F_M.MRAM[799][3] ),
    .B(_2130_),
    .ZN(_2131_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5486_ (.A1(_1799_),
    .A2(_2075_),
    .ZN(_2132_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5487_ (.A1(_2072_),
    .A2(_2132_),
    .ZN(_2133_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _5488_ (.A1(_2114_),
    .A2(_2128_),
    .B1(_2131_),
    .B2(_2133_),
    .ZN(_0035_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5489_ (.I(_2059_),
    .Z(_2134_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5490_ (.I(_2134_),
    .Z(_2135_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _5491_ (.A1(_1791_),
    .A2(\mod.Data_Mem.F_M.MRAM[31][4] ),
    .Z(_2136_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _5492_ (.A1(_2135_),
    .A2(\mod.Data_Mem.F_M.MRAM[30][4] ),
    .B(_2136_),
    .ZN(_2137_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _5493_ (.I(_1690_),
    .Z(_2138_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _5494_ (.A1(_1677_),
    .A2(\mod.Data_Mem.F_M.MRAM[799][4] ),
    .Z(_2139_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _5495_ (.A1(_2138_),
    .A2(\mod.Data_Mem.F_M.MRAM[798][4] ),
    .B(_2139_),
    .ZN(_2140_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _5496_ (.A1(_2119_),
    .A2(_2137_),
    .B1(_2140_),
    .B2(_2133_),
    .ZN(_0036_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _5497_ (.A1(_1686_),
    .A2(\mod.Data_Mem.F_M.MRAM[799][5] ),
    .Z(_2141_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _5498_ (.A1(_1778_),
    .A2(\mod.Data_Mem.F_M.MRAM[798][5] ),
    .B(_2141_),
    .ZN(_2142_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _5499_ (.A1(_1879_),
    .A2(\mod.Data_Mem.F_M.MRAM[30][5] ),
    .Z(_2143_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5500_ (.I(_2059_),
    .Z(_2144_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _5501_ (.A1(_2144_),
    .A2(\mod.Data_Mem.F_M.MRAM[31][5] ),
    .Z(_2145_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5502_ (.A1(_2143_),
    .A2(_2145_),
    .B(_2084_),
    .ZN(_2146_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _5503_ (.A1(_2085_),
    .A2(_2142_),
    .B(_2146_),
    .C(_2104_),
    .ZN(_0037_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _5504_ (.A1(_1791_),
    .A2(\mod.Data_Mem.F_M.MRAM[31][6] ),
    .Z(_2147_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _5505_ (.A1(_2135_),
    .A2(\mod.Data_Mem.F_M.MRAM[30][6] ),
    .B(_2147_),
    .ZN(_2148_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _5506_ (.A1(_1677_),
    .A2(\mod.Data_Mem.F_M.MRAM[799][6] ),
    .Z(_2149_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _5507_ (.A1(_2138_),
    .A2(\mod.Data_Mem.F_M.MRAM[798][6] ),
    .B(_2149_),
    .ZN(_2150_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _5508_ (.A1(_2119_),
    .A2(_2148_),
    .B1(_2150_),
    .B2(_2133_),
    .ZN(_0038_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5509_ (.I(_2144_),
    .Z(_2151_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _5510_ (.I(_1779_),
    .Z(_2152_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _5511_ (.A1(_2152_),
    .A2(\mod.Data_Mem.F_M.MRAM[31][7] ),
    .Z(_2153_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _5512_ (.A1(_2151_),
    .A2(\mod.Data_Mem.F_M.MRAM[30][7] ),
    .B(_2153_),
    .ZN(_2154_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _5513_ (.A1(_1715_),
    .A2(\mod.Data_Mem.F_M.MRAM[799][7] ),
    .Z(_2155_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _5514_ (.A1(_2138_),
    .A2(\mod.Data_Mem.F_M.MRAM[798][7] ),
    .B(_2155_),
    .ZN(_2156_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _5515_ (.A1(_2119_),
    .A2(_2154_),
    .B1(_2156_),
    .B2(_2133_),
    .ZN(_0039_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5516_ (.I(_1543_),
    .Z(_2157_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5517_ (.I(_2157_),
    .Z(_2158_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5518_ (.A1(_2158_),
    .A2(_2093_),
    .ZN(_2159_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5519_ (.I(_1527_),
    .Z(_2160_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _5520_ (.I(_1942_),
    .Z(_2161_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5521_ (.I(_1812_),
    .Z(_2162_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5522_ (.A1(_2161_),
    .A2(\mod.Data_Mem.F_M.MRAM[30][0] ),
    .B1(\mod.Data_Mem.F_M.MRAM[31][0] ),
    .B2(_2162_),
    .ZN(_2163_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5523_ (.I(_2163_),
    .ZN(_2164_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5524_ (.A1(\mod.Data_Mem.F_M.MRAM[29][0] ),
    .A2(_2087_),
    .B1(_2160_),
    .B2(_2164_),
    .ZN(_2165_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5525_ (.I(_2114_),
    .ZN(_2166_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _5526_ (.A1(_2081_),
    .A2(_2067_),
    .B1(_2159_),
    .B2(_2165_),
    .C(_2166_),
    .ZN(_2167_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5527_ (.I(_2132_),
    .Z(_2168_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5528_ (.I(_1713_),
    .Z(_2169_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5529_ (.I(_1915_),
    .Z(_2170_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5530_ (.I(_1782_),
    .Z(_2171_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _5531_ (.A1(_2170_),
    .A2(\mod.Data_Mem.F_M.MRAM[798][0] ),
    .B1(\mod.Data_Mem.F_M.MRAM[799][0] ),
    .B2(_2171_),
    .ZN(_2172_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5532_ (.A1(_2169_),
    .A2(_2172_),
    .ZN(_2173_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5533_ (.A1(\mod.Data_Mem.F_M.MRAM[797][0] ),
    .A2(_1729_),
    .B(_2173_),
    .ZN(_2174_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _5534_ (.A1(_2158_),
    .A2(_2168_),
    .A3(_2174_),
    .ZN(_2175_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _5535_ (.A1(_2167_),
    .A2(_2175_),
    .Z(_2176_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5536_ (.I(_2176_),
    .Z(_0040_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5537_ (.A1(_2158_),
    .A2(_2132_),
    .ZN(_2177_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5538_ (.I(_2177_),
    .Z(_2178_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _5539_ (.I(_2086_),
    .Z(_2179_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5540_ (.I(_1572_),
    .Z(_2180_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _5541_ (.A1(_1782_),
    .A2(\mod.Data_Mem.F_M.MRAM[799][1] ),
    .B1(\mod.Data_Mem.F_M.MRAM[798][1] ),
    .B2(_2009_),
    .ZN(_2181_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5542_ (.A1(_2180_),
    .A2(_2181_),
    .ZN(_2182_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _5543_ (.A1(\mod.Data_Mem.F_M.MRAM[797][1] ),
    .A2(_2179_),
    .B1(_1640_),
    .B2(\mod.Data_Mem.F_M.MRAM[796][1] ),
    .C(_2182_),
    .ZN(_2183_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5544_ (.I(_1804_),
    .Z(_2184_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5545_ (.I(_1533_),
    .Z(_2185_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5546_ (.I(_1602_),
    .Z(_2186_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5547_ (.I(_1914_),
    .Z(_2187_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5548_ (.I(_2187_),
    .Z(_2188_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5549_ (.I(_1790_),
    .Z(_2189_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _5550_ (.A1(_2188_),
    .A2(\mod.Data_Mem.F_M.MRAM[30][1] ),
    .B1(_1632_),
    .B2(_2189_),
    .ZN(_2190_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5551_ (.A1(_2186_),
    .A2(_2190_),
    .ZN(_2191_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_2 _5552_ (.A1(\mod.Data_Mem.F_M.MRAM[29][1] ),
    .A2(_1539_),
    .B1(_1809_),
    .B2(\mod.Data_Mem.F_M.MRAM[28][1] ),
    .C(_2191_),
    .ZN(_2192_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _5553_ (.A1(_2169_),
    .A2(_2185_),
    .B1(_2159_),
    .B2(_2192_),
    .ZN(_2193_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5554_ (.A1(_2184_),
    .A2(_2193_),
    .ZN(_2194_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5555_ (.A1(_2178_),
    .A2(_2183_),
    .B(_2194_),
    .ZN(_0041_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _5556_ (.I(_1639_),
    .Z(_2195_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5557_ (.I(_1644_),
    .Z(_2196_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _5558_ (.A1(_2189_),
    .A2(\mod.Data_Mem.F_M.MRAM[799][2] ),
    .B1(\mod.Data_Mem.F_M.MRAM[798][2] ),
    .B2(_1915_),
    .ZN(_2197_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5559_ (.A1(_2196_),
    .A2(_2197_),
    .ZN(_2198_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _5560_ (.A1(\mod.Data_Mem.F_M.MRAM[797][2] ),
    .A2(_2179_),
    .B1(_2195_),
    .B2(\mod.Data_Mem.F_M.MRAM[796][2] ),
    .C(_2198_),
    .ZN(_2199_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5561_ (.I(_1538_),
    .Z(_2200_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5562_ (.I(_1542_),
    .Z(_2201_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5563_ (.I(_2201_),
    .Z(_2202_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5564_ (.I(_2096_),
    .Z(_2203_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5565_ (.A1(_2070_),
    .A2(\mod.Data_Mem.F_M.MRAM[30][2] ),
    .B1(\mod.Data_Mem.F_M.MRAM[31][2] ),
    .B2(_2203_),
    .ZN(_2204_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5566_ (.A1(_1664_),
    .A2(_2204_),
    .ZN(_2205_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_2 _5567_ (.A1(\mod.Data_Mem.F_M.MRAM[29][2] ),
    .A2(_2200_),
    .B1(_2202_),
    .B2(\mod.Data_Mem.F_M.MRAM[28][2] ),
    .C(_2205_),
    .ZN(_2206_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5568_ (.A1(_2159_),
    .A2(_2206_),
    .B(_1631_),
    .ZN(_2207_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5569_ (.A1(_2184_),
    .A2(_2207_),
    .ZN(_2208_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5570_ (.A1(_2178_),
    .A2(_2199_),
    .B(_2208_),
    .ZN(_0042_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5571_ (.I(_1548_),
    .Z(_2209_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5572_ (.I(_2209_),
    .Z(_2210_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5573_ (.I(_2210_),
    .Z(_2211_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5574_ (.I(_1601_),
    .Z(_2212_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5575_ (.I(\mod.Data_Mem.F_M.MRAM[29][3] ),
    .ZN(_2213_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5576_ (.I(_2060_),
    .Z(_2214_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5577_ (.A1(_2214_),
    .A2(\mod.Data_Mem.F_M.MRAM[31][3] ),
    .ZN(_2215_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5578_ (.I(_1493_),
    .Z(_2216_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5579_ (.I(_2216_),
    .Z(_2217_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5580_ (.A1(_2061_),
    .A2(\mod.Data_Mem.F_M.MRAM[30][3] ),
    .B(_2217_),
    .ZN(_2218_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5581_ (.A1(_2213_),
    .A2(_2179_),
    .B1(_2215_),
    .B2(_2218_),
    .ZN(_2219_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _5582_ (.A1(_2211_),
    .A2(_2212_),
    .A3(_2219_),
    .ZN(_2220_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5583_ (.I(_1549_),
    .Z(_2221_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5584_ (.A1(_2138_),
    .A2(\mod.Data_Mem.F_M.MRAM[799][3] ),
    .B1(\mod.Data_Mem.F_M.MRAM[798][3] ),
    .B2(_2088_),
    .ZN(_2222_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5585_ (.A1(_2221_),
    .A2(_2222_),
    .ZN(_2223_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _5586_ (.A1(\mod.Data_Mem.F_M.MRAM[797][3] ),
    .A2(_2179_),
    .B1(_2195_),
    .B2(\mod.Data_Mem.F_M.MRAM[796][3] ),
    .C(_2223_),
    .ZN(_2224_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _5587_ (.A1(_2114_),
    .A2(_2220_),
    .B1(_2224_),
    .B2(_2178_),
    .ZN(_0043_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _5588_ (.A1(_1800_),
    .A2(_2158_),
    .A3(_2093_),
    .ZN(_2225_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _5589_ (.I(_1549_),
    .Z(_2226_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _5590_ (.I(_1600_),
    .Z(_2227_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5591_ (.I(_1606_),
    .Z(_2228_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5592_ (.I(_1811_),
    .Z(_2229_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _5593_ (.A1(_1953_),
    .A2(\mod.Data_Mem.F_M.MRAM[31][4] ),
    .B1(\mod.Data_Mem.F_M.MRAM[30][4] ),
    .B2(_2229_),
    .ZN(_2230_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5594_ (.A1(_2228_),
    .A2(_2230_),
    .ZN(_2231_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _5595_ (.A1(\mod.Data_Mem.F_M.MRAM[29][4] ),
    .A2(_2226_),
    .B1(_2227_),
    .B2(\mod.Data_Mem.F_M.MRAM[28][4] ),
    .C(_2231_),
    .ZN(_2232_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5596_ (.I(_1594_),
    .Z(_2233_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5597_ (.I(_1811_),
    .Z(_2234_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _5598_ (.A1(_2233_),
    .A2(\mod.Data_Mem.F_M.MRAM[799][4] ),
    .B1(\mod.Data_Mem.F_M.MRAM[798][4] ),
    .B2(_2234_),
    .ZN(_2235_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5599_ (.A1(_1574_),
    .A2(_2235_),
    .ZN(_2236_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _5600_ (.A1(\mod.Data_Mem.F_M.MRAM[797][4] ),
    .A2(_2221_),
    .B1(_1749_),
    .B2(\mod.Data_Mem.F_M.MRAM[796][4] ),
    .C(_2236_),
    .ZN(_2237_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _5601_ (.A1(_2225_),
    .A2(_2232_),
    .B1(_2237_),
    .B2(_2178_),
    .ZN(_0044_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _5602_ (.A1(_1953_),
    .A2(\mod.Data_Mem.F_M.MRAM[31][5] ),
    .B1(\mod.Data_Mem.F_M.MRAM[30][5] ),
    .B2(_2229_),
    .ZN(_2238_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5603_ (.A1(_2228_),
    .A2(_2238_),
    .ZN(_2239_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _5604_ (.A1(\mod.Data_Mem.F_M.MRAM[29][5] ),
    .A2(_2226_),
    .B1(_2227_),
    .B2(\mod.Data_Mem.F_M.MRAM[28][5] ),
    .C(_2239_),
    .ZN(_2240_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _5605_ (.A1(_2233_),
    .A2(\mod.Data_Mem.F_M.MRAM[799][5] ),
    .B1(\mod.Data_Mem.F_M.MRAM[798][5] ),
    .B2(_2234_),
    .ZN(_2241_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5606_ (.A1(_1940_),
    .A2(_2241_),
    .ZN(_2242_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _5607_ (.A1(\mod.Data_Mem.F_M.MRAM[797][5] ),
    .A2(_2221_),
    .B1(_1749_),
    .B2(\mod.Data_Mem.F_M.MRAM[796][5] ),
    .C(_2242_),
    .ZN(_2243_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _5608_ (.A1(_2225_),
    .A2(_2240_),
    .B1(_2243_),
    .B2(_2177_),
    .ZN(_0045_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _5609_ (.A1(_1953_),
    .A2(\mod.Data_Mem.F_M.MRAM[31][6] ),
    .B1(\mod.Data_Mem.F_M.MRAM[30][6] ),
    .B2(_2229_),
    .ZN(_2244_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5610_ (.A1(_2228_),
    .A2(_2244_),
    .ZN(_2245_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _5611_ (.A1(\mod.Data_Mem.F_M.MRAM[29][6] ),
    .A2(_2086_),
    .B1(_2227_),
    .B2(\mod.Data_Mem.F_M.MRAM[28][6] ),
    .C(_2245_),
    .ZN(_2246_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _5612_ (.A1(_2233_),
    .A2(\mod.Data_Mem.F_M.MRAM[799][6] ),
    .B1(\mod.Data_Mem.F_M.MRAM[798][6] ),
    .B2(_2234_),
    .ZN(_2247_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5613_ (.A1(_1940_),
    .A2(_2247_),
    .ZN(_2248_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _5614_ (.A1(\mod.Data_Mem.F_M.MRAM[797][6] ),
    .A2(_2226_),
    .B1(_1749_),
    .B2(\mod.Data_Mem.F_M.MRAM[796][6] ),
    .C(_2248_),
    .ZN(_2249_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _5615_ (.A1(_2225_),
    .A2(_2246_),
    .B1(_2249_),
    .B2(_2177_),
    .ZN(_0046_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _5616_ (.A1(_1746_),
    .A2(\mod.Data_Mem.F_M.MRAM[31][7] ),
    .B1(\mod.Data_Mem.F_M.MRAM[30][7] ),
    .B2(_2187_),
    .ZN(_2250_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5617_ (.A1(_1737_),
    .A2(_2250_),
    .ZN(_2251_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _5618_ (.A1(\mod.Data_Mem.F_M.MRAM[29][7] ),
    .A2(_2086_),
    .B1(_1639_),
    .B2(\mod.Data_Mem.F_M.MRAM[28][7] ),
    .C(_2251_),
    .ZN(_2252_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _5619_ (.A1(_2233_),
    .A2(\mod.Data_Mem.F_M.MRAM[799][7] ),
    .B1(\mod.Data_Mem.F_M.MRAM[798][7] ),
    .B2(_2229_),
    .ZN(_2253_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5620_ (.A1(_1940_),
    .A2(_2253_),
    .ZN(_2254_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _5621_ (.A1(\mod.Data_Mem.F_M.MRAM[797][7] ),
    .A2(_2226_),
    .B1(_2227_),
    .B2(\mod.Data_Mem.F_M.MRAM[796][7] ),
    .C(_2254_),
    .ZN(_2255_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _5622_ (.A1(_2225_),
    .A2(_2252_),
    .B1(_2255_),
    .B2(_2177_),
    .ZN(_0047_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5623_ (.I(_2060_),
    .Z(_2256_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5624_ (.A1(_2256_),
    .A2(\mod.Data_Mem.F_M.MRAM[797][0] ),
    .ZN(_2257_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _5625_ (.I(_1845_),
    .Z(_2258_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5626_ (.I(_2216_),
    .Z(_2259_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5627_ (.A1(_2258_),
    .A2(\mod.Data_Mem.F_M.MRAM[796][0] ),
    .B(_2259_),
    .ZN(_2260_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _5628_ (.A1(_2089_),
    .A2(_2099_),
    .B1(_2257_),
    .B2(_2260_),
    .ZN(_2261_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5629_ (.A1(_2094_),
    .A2(_2261_),
    .ZN(_2262_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5630_ (.I(_2075_),
    .Z(_2263_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5631_ (.I(_1840_),
    .Z(_2264_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5632_ (.A1(_2264_),
    .A2(\mod.Data_Mem.F_M.MRAM[29][0] ),
    .ZN(_2265_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5633_ (.I(_1875_),
    .Z(_2266_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5634_ (.I(_1493_),
    .Z(_2267_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5635_ (.I(_2267_),
    .Z(_2268_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5636_ (.A1(_2266_),
    .A2(\mod.Data_Mem.F_M.MRAM[28][0] ),
    .B(_2268_),
    .ZN(_2269_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5637_ (.I(_1811_),
    .Z(_2270_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5638_ (.A1(_2270_),
    .A2(_2112_),
    .ZN(_2271_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5639_ (.A1(_2265_),
    .A2(_2269_),
    .B(_2271_),
    .ZN(_2272_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _5640_ (.A1(_2084_),
    .A2(_2263_),
    .A3(_2272_),
    .ZN(_2273_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _5641_ (.A1(_2063_),
    .A2(_2113_),
    .B(_2262_),
    .C(_2273_),
    .ZN(_0048_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5642_ (.A1(_2264_),
    .A2(\mod.Data_Mem.F_M.MRAM[797][1] ),
    .ZN(_2274_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5643_ (.I(_1586_),
    .Z(_2275_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5644_ (.A1(_2275_),
    .A2(\mod.Data_Mem.F_M.MRAM[796][1] ),
    .B(_2268_),
    .ZN(_2276_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5645_ (.A1(_2270_),
    .A2(_2122_),
    .ZN(_2277_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5646_ (.A1(_2274_),
    .A2(_2276_),
    .B(_2277_),
    .ZN(_2278_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5647_ (.A1(_2168_),
    .A2(_2278_),
    .ZN(_2279_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5648_ (.I(_2088_),
    .Z(_2280_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5649_ (.I(_2060_),
    .Z(_2281_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5650_ (.A1(_2281_),
    .A2(\mod.Data_Mem.F_M.MRAM[29][1] ),
    .ZN(_2282_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5651_ (.I(_1779_),
    .Z(_2283_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5652_ (.A1(_2283_),
    .A2(\mod.Data_Mem.F_M.MRAM[28][1] ),
    .B(_2217_),
    .ZN(_2284_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _5653_ (.A1(_2280_),
    .A2(_2121_),
    .B1(_2282_),
    .B2(_2284_),
    .ZN(_2285_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5654_ (.A1(_2068_),
    .A2(_2285_),
    .ZN(_2286_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _5655_ (.A1(_2091_),
    .A2(_1803_),
    .B(_2279_),
    .C(_2286_),
    .ZN(_0049_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5656_ (.A1(_2151_),
    .A2(\mod.Data_Mem.F_M.MRAM[797][2] ),
    .ZN(_2287_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5657_ (.I(_1609_),
    .Z(_2288_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5658_ (.A1(_2288_),
    .A2(\mod.Data_Mem.F_M.MRAM[796][2] ),
    .B(_2268_),
    .ZN(_2289_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5659_ (.I(_1914_),
    .Z(_2290_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5660_ (.A1(_2290_),
    .A2(_2125_),
    .ZN(_2291_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5661_ (.A1(_2287_),
    .A2(_2289_),
    .B(_2291_),
    .ZN(_2292_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5662_ (.A1(_2168_),
    .A2(_2292_),
    .ZN(_2293_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5663_ (.A1(_2135_),
    .A2(\mod.Data_Mem.F_M.MRAM[29][2] ),
    .ZN(_2294_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5664_ (.I(_1686_),
    .Z(_2295_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5665_ (.A1(_2295_),
    .A2(\mod.Data_Mem.F_M.MRAM[28][2] ),
    .B(_2259_),
    .ZN(_2296_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5666_ (.A1(_2290_),
    .A2(_2124_),
    .ZN(_2297_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5667_ (.A1(_2294_),
    .A2(_2296_),
    .B(_2297_),
    .ZN(_2298_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5668_ (.A1(_2068_),
    .A2(_2298_),
    .ZN(_2299_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _5669_ (.A1(_2074_),
    .A2(_2118_),
    .B(_2293_),
    .C(_2299_),
    .ZN(_0050_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5670_ (.A1(_2270_),
    .A2(_2127_),
    .ZN(_2300_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5671_ (.I(_1692_),
    .Z(_2301_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5672_ (.A1(_2301_),
    .A2(_2213_),
    .ZN(_2302_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _5673_ (.A1(_2288_),
    .A2(\mod.Data_Mem.F_M.MRAM[28][3] ),
    .B(_2302_),
    .C(_2268_),
    .ZN(_2303_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5674_ (.A1(_2300_),
    .A2(_2303_),
    .ZN(_2304_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5675_ (.A1(_2076_),
    .A2(_2304_),
    .B(_2166_),
    .ZN(_2305_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5676_ (.I(_2132_),
    .Z(_2306_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5677_ (.A1(_2135_),
    .A2(\mod.Data_Mem.F_M.MRAM[797][3] ),
    .ZN(_2307_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5678_ (.A1(_2295_),
    .A2(\mod.Data_Mem.F_M.MRAM[796][3] ),
    .B(_2259_),
    .ZN(_2308_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _5679_ (.A1(_2089_),
    .A2(_2131_),
    .B1(_2307_),
    .B2(_2308_),
    .ZN(_2309_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5680_ (.A1(_2306_),
    .A2(_2309_),
    .ZN(_2310_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5681_ (.A1(_2305_),
    .A2(_2310_),
    .ZN(_0051_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5682_ (.I(_2069_),
    .Z(_2311_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5683_ (.I(_2311_),
    .Z(_2312_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5684_ (.I(_1691_),
    .Z(_2313_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5685_ (.A1(_2313_),
    .A2(\mod.Data_Mem.F_M.MRAM[29][4] ),
    .ZN(_2314_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5686_ (.I(_1675_),
    .Z(_2315_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5687_ (.I(_2267_),
    .Z(_2316_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5688_ (.A1(_2315_),
    .A2(\mod.Data_Mem.F_M.MRAM[28][4] ),
    .B(_2316_),
    .ZN(_2317_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _5689_ (.A1(_2312_),
    .A2(_2137_),
    .B1(_2314_),
    .B2(_2317_),
    .ZN(_2318_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5690_ (.I(_2096_),
    .Z(_2319_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5691_ (.A1(_2319_),
    .A2(\mod.Data_Mem.F_M.MRAM[797][4] ),
    .ZN(_2320_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5692_ (.I(_1593_),
    .Z(_2321_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5693_ (.A1(_2321_),
    .A2(\mod.Data_Mem.F_M.MRAM[796][4] ),
    .B(_2311_),
    .ZN(_2322_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _5694_ (.A1(_2280_),
    .A2(_2140_),
    .B1(_2320_),
    .B2(_2322_),
    .ZN(_2323_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5695_ (.A1(_2082_),
    .A2(_2318_),
    .B1(_2323_),
    .B2(_2306_),
    .ZN(_2324_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5696_ (.I(_2324_),
    .ZN(_0052_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5697_ (.A1(_2256_),
    .A2(\mod.Data_Mem.F_M.MRAM[29][5] ),
    .ZN(_2325_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _5698_ (.I(_1517_),
    .Z(_2326_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5699_ (.A1(_2326_),
    .A2(\mod.Data_Mem.F_M.MRAM[28][5] ),
    .B(_2259_),
    .ZN(_2327_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _5700_ (.A1(_2116_),
    .A2(_2143_),
    .A3(_2145_),
    .ZN(_2328_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5701_ (.A1(_2325_),
    .A2(_2327_),
    .B(_2328_),
    .ZN(_2329_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5702_ (.A1(_2203_),
    .A2(\mod.Data_Mem.F_M.MRAM[797][5] ),
    .ZN(_2330_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _5703_ (.I(_1581_),
    .Z(_2331_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5704_ (.A1(_2331_),
    .A2(\mod.Data_Mem.F_M.MRAM[796][5] ),
    .B(_2088_),
    .ZN(_2332_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _5705_ (.A1(_2316_),
    .A2(_2142_),
    .B1(_2330_),
    .B2(_2332_),
    .ZN(_2333_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5706_ (.A1(_2082_),
    .A2(_2329_),
    .B1(_2333_),
    .B2(_2306_),
    .ZN(_2334_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5707_ (.I(_2334_),
    .ZN(_0053_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5708_ (.A1(_2313_),
    .A2(\mod.Data_Mem.F_M.MRAM[29][6] ),
    .ZN(_2335_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5709_ (.A1(_2315_),
    .A2(\mod.Data_Mem.F_M.MRAM[28][6] ),
    .B(_2316_),
    .ZN(_2336_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _5710_ (.A1(_2071_),
    .A2(_2148_),
    .B1(_2335_),
    .B2(_2336_),
    .ZN(_2337_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5711_ (.A1(_2129_),
    .A2(\mod.Data_Mem.F_M.MRAM[797][6] ),
    .ZN(_2338_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _5712_ (.I(_2025_),
    .Z(_2339_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5713_ (.A1(_2339_),
    .A2(\mod.Data_Mem.F_M.MRAM[796][6] ),
    .B(_2311_),
    .ZN(_2340_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _5714_ (.A1(_2316_),
    .A2(_2150_),
    .B1(_2338_),
    .B2(_2340_),
    .ZN(_2341_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5715_ (.A1(_2082_),
    .A2(_2337_),
    .B1(_2341_),
    .B2(_2306_),
    .ZN(_2342_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5716_ (.I(_2342_),
    .ZN(_0054_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5717_ (.I(_1691_),
    .Z(_2343_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5718_ (.A1(_2343_),
    .A2(\mod.Data_Mem.F_M.MRAM[29][7] ),
    .ZN(_2344_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5719_ (.I(_1714_),
    .Z(_2345_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5720_ (.A1(_2345_),
    .A2(\mod.Data_Mem.F_M.MRAM[28][7] ),
    .B(_2280_),
    .ZN(_2346_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _5721_ (.A1(_2312_),
    .A2(_2154_),
    .B1(_2344_),
    .B2(_2346_),
    .ZN(_2347_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5722_ (.A1(_2281_),
    .A2(\mod.Data_Mem.F_M.MRAM[797][7] ),
    .ZN(_2348_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5723_ (.A1(_1932_),
    .A2(\mod.Data_Mem.F_M.MRAM[796][7] ),
    .B(_2217_),
    .ZN(_2349_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _5724_ (.A1(_2280_),
    .A2(_2156_),
    .B1(_2348_),
    .B2(_2349_),
    .ZN(_2350_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5725_ (.A1(_2068_),
    .A2(_2347_),
    .B1(_2350_),
    .B2(_2168_),
    .ZN(_2351_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5726_ (.I(_2351_),
    .ZN(_0055_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5727_ (.I(_2209_),
    .Z(_2352_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5728_ (.I(_2352_),
    .Z(_2353_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5729_ (.A1(_1812_),
    .A2(_1553_),
    .ZN(_2354_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5730_ (.I(_2354_),
    .Z(_2355_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5731_ (.A1(_2187_),
    .A2(_1499_),
    .ZN(_2356_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5732_ (.I(_2356_),
    .Z(_2357_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _5733_ (.I(_1681_),
    .Z(_2358_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5734_ (.I0(\mod.Data_Mem.F_M.MRAM[14][0] ),
    .I1(\mod.Data_Mem.F_M.MRAM[15][0] ),
    .S(_2358_),
    .Z(_2359_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _5735_ (.I(_1677_),
    .Z(_2360_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5736_ (.I0(\mod.Data_Mem.F_M.MRAM[16][0] ),
    .I1(\mod.Data_Mem.F_M.MRAM[17][0] ),
    .S(_2360_),
    .Z(_2361_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5737_ (.I(_2162_),
    .Z(_2362_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _5738_ (.A1(_2112_),
    .A2(_2355_),
    .B1(_2357_),
    .B2(_2359_),
    .C1(_2361_),
    .C2(_2362_),
    .ZN(_2363_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _5739_ (.I0(\mod.Data_Mem.F_M.MRAM[4][0] ),
    .I1(\mod.Data_Mem.F_M.MRAM[5][0] ),
    .I2(\mod.Data_Mem.F_M.MRAM[20][0] ),
    .I3(\mod.Data_Mem.F_M.MRAM[21][0] ),
    .S0(_1714_),
    .S1(_1756_),
    .Z(_2364_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5740_ (.I0(\mod.Data_Mem.F_M.MRAM[18][0] ),
    .I1(\mod.Data_Mem.F_M.MRAM[19][0] ),
    .S(_2358_),
    .Z(_2365_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5741_ (.I(_2064_),
    .Z(_2366_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5742_ (.I(_2356_),
    .Z(_2367_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5743_ (.I0(\mod.Data_Mem.F_M.MRAM[2][0] ),
    .I1(\mod.Data_Mem.F_M.MRAM[3][0] ),
    .S(_1515_),
    .Z(_2368_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5744_ (.A1(_2367_),
    .A2(_2368_),
    .ZN(_2369_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5745_ (.A1(_2366_),
    .A2(_2369_),
    .ZN(_2370_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _5746_ (.A1(_2362_),
    .A2(_2364_),
    .B1(_2365_),
    .B2(_2355_),
    .C(_2370_),
    .ZN(_2371_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _5747_ (.A1(_2353_),
    .A2(_2363_),
    .B(_2371_),
    .C(_1498_),
    .ZN(_2372_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5748_ (.A1(_1542_),
    .A2(_1533_),
    .ZN(_2373_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5749_ (.I(_2373_),
    .Z(_2374_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5750_ (.A1(_1595_),
    .A2(_1500_),
    .ZN(_2375_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5751_ (.I(_2375_),
    .Z(_2376_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5752_ (.A1(_2106_),
    .A2(_2376_),
    .ZN(_2377_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5753_ (.I(_2377_),
    .Z(_2378_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5754_ (.I(_2378_),
    .Z(_2379_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5755_ (.A1(_2187_),
    .A2(_2064_),
    .ZN(_2380_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5756_ (.I(_2380_),
    .Z(_2381_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5757_ (.I(_2381_),
    .Z(_2382_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5758_ (.I(_1588_),
    .Z(_2383_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5759_ (.I0(\mod.Data_Mem.F_M.MRAM[782][0] ),
    .I1(\mod.Data_Mem.F_M.MRAM[783][0] ),
    .S(_2383_),
    .Z(_2384_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5760_ (.I(_1840_),
    .Z(_2385_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _5761_ (.A1(_1954_),
    .A2(\mod.Data_Mem.F_M.MRAM[769][0] ),
    .Z(_2386_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5762_ (.A1(_2385_),
    .A2(\mod.Data_Mem.F_M.MRAM[768][0] ),
    .B(_2386_),
    .ZN(_2387_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5763_ (.I(_2101_),
    .Z(_2388_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5764_ (.I0(\mod.Data_Mem.F_M.MRAM[770][0] ),
    .I1(\mod.Data_Mem.F_M.MRAM[771][0] ),
    .S(_1581_),
    .Z(_2389_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5765_ (.I0(\mod.Data_Mem.F_M.MRAM[772][0] ),
    .I1(\mod.Data_Mem.F_M.MRAM[773][0] ),
    .S(_1951_),
    .Z(_2390_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _5766_ (.A1(_2388_),
    .A2(_2389_),
    .B1(_2390_),
    .B2(_2290_),
    .C(_2376_),
    .ZN(_2391_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5767_ (.A1(_2210_),
    .A2(_2387_),
    .B(_2391_),
    .ZN(_2392_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5768_ (.A1(_2382_),
    .A2(_2384_),
    .B(_2392_),
    .ZN(_2393_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5769_ (.I(_2380_),
    .Z(_2394_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5770_ (.A1(_1595_),
    .A2(_1554_),
    .ZN(_2395_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5771_ (.I(_2395_),
    .Z(_2396_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5772_ (.I(_2396_),
    .Z(_2397_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _5773_ (.I(_1658_),
    .Z(_2398_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _5774_ (.A1(_2398_),
    .A2(\mod.Data_Mem.F_M.MRAM[789][0] ),
    .Z(_2399_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5775_ (.A1(_2313_),
    .A2(\mod.Data_Mem.F_M.MRAM[788][0] ),
    .B(_2399_),
    .ZN(_2400_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5776_ (.A1(_2394_),
    .A2(_2099_),
    .B1(_2397_),
    .B2(_2400_),
    .ZN(_2401_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5777_ (.A1(_2008_),
    .A2(_1548_),
    .ZN(_2402_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5778_ (.I(_2402_),
    .Z(_2403_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5779_ (.I0(\mod.Data_Mem.F_M.MRAM[784][0] ),
    .I1(\mod.Data_Mem.F_M.MRAM[785][0] ),
    .S(_1791_),
    .Z(_2404_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5780_ (.A1(_2403_),
    .A2(_2404_),
    .ZN(_2405_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5781_ (.I(_2109_),
    .Z(_2406_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5782_ (.I0(\mod.Data_Mem.F_M.MRAM[786][0] ),
    .I1(\mod.Data_Mem.F_M.MRAM[787][0] ),
    .S(_1769_),
    .Z(_2407_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5783_ (.A1(_2406_),
    .A2(_2407_),
    .ZN(_2408_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5784_ (.A1(_2405_),
    .A2(_2408_),
    .ZN(_2409_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5785_ (.I(_2377_),
    .Z(_2410_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5786_ (.A1(_2401_),
    .A2(_2409_),
    .B(_2410_),
    .ZN(_2411_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5787_ (.A1(_2379_),
    .A2(_2393_),
    .B(_2411_),
    .ZN(_2412_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5788_ (.A1(_1490_),
    .A2(_2117_),
    .ZN(_2413_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5789_ (.I(_2413_),
    .Z(_2414_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _5790_ (.A1(_1491_),
    .A2(_2372_),
    .A3(_2374_),
    .B1(_2412_),
    .B2(_2414_),
    .ZN(_2415_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5791_ (.I(_2415_),
    .ZN(_0056_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5792_ (.I(_2378_),
    .Z(_2416_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5793_ (.I(_1675_),
    .Z(_2417_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5794_ (.I(_1517_),
    .Z(_2418_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5795_ (.A1(_2418_),
    .A2(\mod.Data_Mem.F_M.MRAM[787][1] ),
    .ZN(_2419_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5796_ (.A1(_2417_),
    .A2(_1682_),
    .B(_2419_),
    .ZN(_2420_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5797_ (.A1(_2110_),
    .A2(_2420_),
    .ZN(_2421_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5798_ (.I(_1596_),
    .Z(_2422_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5799_ (.I(_2422_),
    .Z(_2423_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5800_ (.I(_1612_),
    .Z(_2424_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5801_ (.I(_1636_),
    .Z(_2425_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5802_ (.A1(_2425_),
    .A2(\mod.Data_Mem.F_M.MRAM[785][1] ),
    .ZN(_2426_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5803_ (.A1(_2424_),
    .A2(_1678_),
    .B(_2426_),
    .ZN(_2427_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5804_ (.I(_1903_),
    .Z(_2428_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5805_ (.I(_2395_),
    .Z(_2429_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5806_ (.A1(_2358_),
    .A2(\mod.Data_Mem.F_M.MRAM[789][1] ),
    .ZN(_2430_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _5807_ (.A1(_2428_),
    .A2(_1687_),
    .B(_2429_),
    .C(_2430_),
    .ZN(_2431_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _5808_ (.A1(_2423_),
    .A2(_2122_),
    .B1(_2427_),
    .B2(_2403_),
    .C(_2431_),
    .ZN(_2432_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5809_ (.A1(_2421_),
    .A2(_2432_),
    .ZN(_2433_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5810_ (.I(_2100_),
    .Z(_2434_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5811_ (.I(_2109_),
    .Z(_2435_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5812_ (.A1(_2152_),
    .A2(\mod.Data_Mem.F_M.MRAM[771][1] ),
    .ZN(_2436_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5813_ (.A1(_2321_),
    .A2(_1709_),
    .B(_2436_),
    .ZN(_2437_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5814_ (.I0(\mod.Data_Mem.F_M.MRAM[782][1] ),
    .I1(\mod.Data_Mem.F_M.MRAM[783][1] ),
    .S(_1918_),
    .Z(_2438_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5815_ (.I(_2422_),
    .Z(_2439_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5816_ (.I(_2396_),
    .Z(_2440_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5817_ (.A1(_2281_),
    .A2(\mod.Data_Mem.F_M.MRAM[772][1] ),
    .ZN(_2441_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5818_ (.A1(_2283_),
    .A2(\mod.Data_Mem.F_M.MRAM[773][1] ),
    .ZN(_2442_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _5819_ (.A1(_2440_),
    .A2(_2441_),
    .A3(_2442_),
    .ZN(_2443_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _5820_ (.A1(_2435_),
    .A2(_2437_),
    .B1(_2438_),
    .B2(_2439_),
    .C(_2443_),
    .ZN(_2444_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5821_ (.A1(_2434_),
    .A2(_2444_),
    .ZN(_2445_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5822_ (.A1(_2416_),
    .A2(_2433_),
    .B(_2445_),
    .ZN(_2446_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5823_ (.I(_2352_),
    .Z(_2447_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _5824_ (.I(_2234_),
    .Z(_2448_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5825_ (.I(_2448_),
    .Z(_2449_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _5826_ (.I0(\mod.Data_Mem.F_M.MRAM[4][1] ),
    .I1(\mod.Data_Mem.F_M.MRAM[5][1] ),
    .I2(\mod.Data_Mem.F_M.MRAM[20][1] ),
    .I3(\mod.Data_Mem.F_M.MRAM[21][1] ),
    .S0(_2025_),
    .S1(_2106_),
    .Z(_2450_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5827_ (.I0(\mod.Data_Mem.F_M.MRAM[2][1] ),
    .I1(\mod.Data_Mem.F_M.MRAM[3][1] ),
    .S(_1954_),
    .Z(_2451_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _5828_ (.I(_1519_),
    .Z(_2452_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5829_ (.I0(\mod.Data_Mem.F_M.MRAM[18][1] ),
    .I1(\mod.Data_Mem.F_M.MRAM[19][1] ),
    .S(_2452_),
    .Z(_2453_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5830_ (.I(_2354_),
    .Z(_2454_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _5831_ (.A1(_2449_),
    .A2(_2450_),
    .B1(_2451_),
    .B2(_2357_),
    .C1(_2453_),
    .C2(_2454_),
    .ZN(_2455_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5832_ (.A1(_2447_),
    .A2(_2455_),
    .ZN(_2456_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5833_ (.I(_2366_),
    .Z(_2457_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5834_ (.I0(\mod.Data_Mem.F_M.MRAM[30][1] ),
    .I1(_1632_),
    .S(_2398_),
    .Z(_2458_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5835_ (.I0(\mod.Data_Mem.F_M.MRAM[14][1] ),
    .I1(\mod.Data_Mem.F_M.MRAM[15][1] ),
    .S(_2452_),
    .Z(_2459_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5836_ (.I0(\mod.Data_Mem.F_M.MRAM[16][1] ),
    .I1(\mod.Data_Mem.F_M.MRAM[17][1] ),
    .S(_2152_),
    .Z(_2460_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _5837_ (.A1(_2458_),
    .A2(_2454_),
    .B1(_2367_),
    .B2(_2459_),
    .C1(_2460_),
    .C2(_2170_),
    .ZN(_2461_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5838_ (.A1(_2457_),
    .A2(_2461_),
    .B(_1804_),
    .ZN(_2462_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5839_ (.A1(_2456_),
    .A2(_2462_),
    .ZN(_2463_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _5840_ (.A1(_2085_),
    .A2(_2446_),
    .B(_2463_),
    .C(_1498_),
    .ZN(_0057_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5841_ (.I(_2109_),
    .Z(_2464_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5842_ (.A1(_2418_),
    .A2(\mod.Data_Mem.F_M.MRAM[787][2] ),
    .ZN(_2465_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5843_ (.A1(_2417_),
    .A2(_1787_),
    .B(_2465_),
    .ZN(_2466_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5844_ (.A1(_2464_),
    .A2(_2466_),
    .ZN(_2467_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5845_ (.A1(_2425_),
    .A2(\mod.Data_Mem.F_M.MRAM[785][2] ),
    .ZN(_2468_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5846_ (.A1(_2424_),
    .A2(_1792_),
    .B(_2468_),
    .ZN(_2469_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5847_ (.A1(_2358_),
    .A2(\mod.Data_Mem.F_M.MRAM[789][2] ),
    .ZN(_2470_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _5848_ (.A1(_2428_),
    .A2(_1784_),
    .B(_2429_),
    .C(_2470_),
    .ZN(_2471_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _5849_ (.A1(_2439_),
    .A2(_2125_),
    .B1(_2469_),
    .B2(_2403_),
    .C(_2471_),
    .ZN(_2472_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5850_ (.A1(_2467_),
    .A2(_2472_),
    .ZN(_2473_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5851_ (.I(_1535_),
    .Z(_2474_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5852_ (.I(_1814_),
    .Z(_2475_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5853_ (.A1(_2161_),
    .A2(\mod.Data_Mem.F_M.MRAM[771][2] ),
    .ZN(_2476_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5854_ (.A1(_2475_),
    .A2(_1765_),
    .B(_2476_),
    .ZN(_2477_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5855_ (.I0(\mod.Data_Mem.F_M.MRAM[782][2] ),
    .I1(\mod.Data_Mem.F_M.MRAM[783][2] ),
    .S(_2398_),
    .Z(_2478_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5856_ (.A1(_2281_),
    .A2(\mod.Data_Mem.F_M.MRAM[772][2] ),
    .ZN(_2479_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5857_ (.A1(_2383_),
    .A2(\mod.Data_Mem.F_M.MRAM[773][2] ),
    .ZN(_2480_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _5858_ (.A1(_2440_),
    .A2(_2479_),
    .A3(_2480_),
    .ZN(_2481_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _5859_ (.A1(_2435_),
    .A2(_2477_),
    .B1(_2478_),
    .B2(_2439_),
    .C(_2481_),
    .ZN(_2482_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5860_ (.A1(_2474_),
    .A2(_2482_),
    .ZN(_2483_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5861_ (.A1(_2416_),
    .A2(_2473_),
    .B(_2483_),
    .ZN(_2484_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _5862_ (.I0(\mod.Data_Mem.F_M.MRAM[4][2] ),
    .I1(\mod.Data_Mem.F_M.MRAM[5][2] ),
    .I2(\mod.Data_Mem.F_M.MRAM[20][2] ),
    .I3(\mod.Data_Mem.F_M.MRAM[21][2] ),
    .S0(_2025_),
    .S1(_2106_),
    .Z(_2485_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5863_ (.I0(\mod.Data_Mem.F_M.MRAM[2][2] ),
    .I1(\mod.Data_Mem.F_M.MRAM[3][2] ),
    .S(_1954_),
    .Z(_2486_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5864_ (.I0(\mod.Data_Mem.F_M.MRAM[18][2] ),
    .I1(\mod.Data_Mem.F_M.MRAM[19][2] ),
    .S(_2452_),
    .Z(_2487_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _5865_ (.A1(_2449_),
    .A2(_2485_),
    .B1(_2486_),
    .B2(_2367_),
    .C1(_2487_),
    .C2(_2454_),
    .ZN(_2488_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5866_ (.A1(_2447_),
    .A2(_2488_),
    .ZN(_2489_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5867_ (.I0(\mod.Data_Mem.F_M.MRAM[14][2] ),
    .I1(\mod.Data_Mem.F_M.MRAM[15][2] ),
    .S(_2452_),
    .Z(_2490_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5868_ (.I0(\mod.Data_Mem.F_M.MRAM[16][2] ),
    .I1(\mod.Data_Mem.F_M.MRAM[17][2] ),
    .S(_2152_),
    .Z(_2491_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _5869_ (.A1(_2124_),
    .A2(_2454_),
    .B1(_2367_),
    .B2(_2490_),
    .C1(_2491_),
    .C2(_2170_),
    .ZN(_2492_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5870_ (.A1(_2457_),
    .A2(_2492_),
    .B(_1804_),
    .ZN(_2493_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5871_ (.A1(_2489_),
    .A2(_2493_),
    .ZN(_2494_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _5872_ (.A1(_2085_),
    .A2(_2484_),
    .B(_2494_),
    .C(_1498_),
    .ZN(_0058_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5873_ (.I(_2101_),
    .Z(_2495_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5874_ (.I(_2495_),
    .Z(_2496_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5875_ (.I0(\mod.Data_Mem.F_M.MRAM[786][3] ),
    .I1(\mod.Data_Mem.F_M.MRAM[787][3] ),
    .S(_1932_),
    .Z(_2497_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5876_ (.A1(_2496_),
    .A2(_2497_),
    .B(_2378_),
    .ZN(_2498_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5877_ (.I(_2395_),
    .Z(_2499_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5878_ (.I(_2499_),
    .Z(_2500_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5879_ (.I0(\mod.Data_Mem.F_M.MRAM[788][3] ),
    .I1(\mod.Data_Mem.F_M.MRAM[789][3] ),
    .S(_2161_),
    .Z(_2501_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5880_ (.I0(\mod.Data_Mem.F_M.MRAM[784][3] ),
    .I1(\mod.Data_Mem.F_M.MRAM[785][3] ),
    .S(_2339_),
    .Z(_2502_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5881_ (.I(_2376_),
    .Z(_2503_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5882_ (.A1(_2500_),
    .A2(_2501_),
    .B1(_2502_),
    .B2(_2503_),
    .ZN(_2504_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _5883_ (.A1(_2423_),
    .A2(_2131_),
    .B(_2498_),
    .C(_2504_),
    .ZN(_2505_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5884_ (.I(_2319_),
    .Z(_2506_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _5885_ (.A1(_2266_),
    .A2(\mod.Data_Mem.F_M.MRAM[782][3] ),
    .Z(_2507_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5886_ (.I(_2209_),
    .Z(_2508_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _5887_ (.A1(_2506_),
    .A2(\mod.Data_Mem.F_M.MRAM[783][3] ),
    .B(_2507_),
    .C(_2508_),
    .ZN(_2509_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5888_ (.I(_2495_),
    .Z(_2510_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5889_ (.I(_1707_),
    .Z(_2511_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5890_ (.I(_1513_),
    .Z(_2512_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5891_ (.A1(_2512_),
    .A2(\mod.Data_Mem.F_M.MRAM[771][3] ),
    .ZN(_2513_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5892_ (.A1(_2511_),
    .A2(_1851_),
    .B(_2513_),
    .ZN(_2514_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5893_ (.A1(_2275_),
    .A2(\mod.Data_Mem.F_M.MRAM[773][3] ),
    .ZN(_2515_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5894_ (.A1(_2511_),
    .A2(_1846_),
    .B(_2515_),
    .ZN(_2516_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5895_ (.I(_2116_),
    .Z(_2517_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5896_ (.A1(_2510_),
    .A2(_2514_),
    .B1(_2516_),
    .B2(_2517_),
    .ZN(_2518_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _5897_ (.A1(_2416_),
    .A2(_2509_),
    .A3(_2518_),
    .ZN(_2519_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _5898_ (.A1(_2118_),
    .A2(_2505_),
    .A3(_2519_),
    .ZN(_2520_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _5899_ (.I0(\mod.Data_Mem.F_M.MRAM[4][3] ),
    .I1(\mod.Data_Mem.F_M.MRAM[5][3] ),
    .I2(\mod.Data_Mem.F_M.MRAM[20][3] ),
    .I3(\mod.Data_Mem.F_M.MRAM[21][3] ),
    .S0(_1918_),
    .S1(_1756_),
    .Z(_2521_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _5900_ (.I(_1609_),
    .Z(_2522_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5901_ (.I0(\mod.Data_Mem.F_M.MRAM[18][3] ),
    .I1(\mod.Data_Mem.F_M.MRAM[19][3] ),
    .S(_2522_),
    .Z(_2523_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5902_ (.I0(\mod.Data_Mem.F_M.MRAM[2][3] ),
    .I1(\mod.Data_Mem.F_M.MRAM[3][3] ),
    .S(_2321_),
    .Z(_2524_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _5903_ (.A1(_2517_),
    .A2(_2521_),
    .B1(_2523_),
    .B2(_2355_),
    .C1(_2524_),
    .C2(_2357_),
    .ZN(_2525_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5904_ (.A1(_2211_),
    .A2(_2525_),
    .ZN(_2526_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5905_ (.I0(\mod.Data_Mem.F_M.MRAM[14][3] ),
    .I1(\mod.Data_Mem.F_M.MRAM[15][3] ),
    .S(_2331_),
    .Z(_2527_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _5906_ (.I(_1894_),
    .Z(_2528_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5907_ (.I0(\mod.Data_Mem.F_M.MRAM[16][3] ),
    .I1(\mod.Data_Mem.F_M.MRAM[17][3] ),
    .S(_2528_),
    .Z(_2529_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _5908_ (.A1(_2127_),
    .A2(_2355_),
    .B1(_2357_),
    .B2(_2527_),
    .C1(_2529_),
    .C2(_2362_),
    .ZN(_2530_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5909_ (.I(_2117_),
    .Z(_2531_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _5910_ (.A1(_2457_),
    .A2(_2530_),
    .B(_2531_),
    .C(_1800_),
    .ZN(_2532_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5911_ (.A1(_2526_),
    .A2(_2532_),
    .ZN(_2533_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5912_ (.A1(_2080_),
    .A2(_2520_),
    .B(_2533_),
    .ZN(_0059_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5913_ (.I(_1726_),
    .Z(_2534_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5914_ (.I(_2394_),
    .Z(_2535_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5915_ (.I(_2440_),
    .Z(_2536_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _5916_ (.A1(_2428_),
    .A2(\mod.Data_Mem.F_M.MRAM[789][4] ),
    .Z(_2537_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5917_ (.A1(_2506_),
    .A2(\mod.Data_Mem.F_M.MRAM[788][4] ),
    .B(_2537_),
    .ZN(_2538_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5918_ (.I(_2402_),
    .Z(_2539_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _5919_ (.I(_1783_),
    .Z(_2540_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5920_ (.I0(\mod.Data_Mem.F_M.MRAM[784][4] ),
    .I1(\mod.Data_Mem.F_M.MRAM[785][4] ),
    .S(_2540_),
    .Z(_2541_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5921_ (.A1(_2097_),
    .A2(\mod.Data_Mem.F_M.MRAM[786][4] ),
    .ZN(_2542_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5922_ (.A1(_2151_),
    .A2(_1919_),
    .B(_2542_),
    .ZN(_2543_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _5923_ (.A1(_2539_),
    .A2(_2541_),
    .B1(_2543_),
    .B2(_2435_),
    .ZN(_2544_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _5924_ (.A1(_2535_),
    .A2(_2140_),
    .B1(_2536_),
    .B2(_2538_),
    .C(_2544_),
    .ZN(_2545_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5925_ (.I0(\mod.Data_Mem.F_M.MRAM[782][4] ),
    .I1(_1901_),
    .S(_2258_),
    .Z(_2546_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5926_ (.I0(\mod.Data_Mem.F_M.MRAM[770][4] ),
    .I1(\mod.Data_Mem.F_M.MRAM[771][4] ),
    .S(_2339_),
    .Z(_2547_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5927_ (.I(_2396_),
    .Z(_2548_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5928_ (.I(_2144_),
    .Z(_2549_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5929_ (.A1(_2549_),
    .A2(\mod.Data_Mem.F_M.MRAM[772][4] ),
    .ZN(_2550_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5930_ (.A1(_2512_),
    .A2(\mod.Data_Mem.F_M.MRAM[773][4] ),
    .ZN(_2551_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _5931_ (.A1(_2548_),
    .A2(_2550_),
    .A3(_2551_),
    .ZN(_2552_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _5932_ (.A1(_2423_),
    .A2(_2546_),
    .B1(_2547_),
    .B2(_2464_),
    .C(_2552_),
    .ZN(_2553_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5933_ (.A1(_2434_),
    .A2(_2553_),
    .ZN(_2554_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5934_ (.A1(_2379_),
    .A2(_2545_),
    .B(_2554_),
    .ZN(_2555_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5935_ (.I0(\mod.Data_Mem.F_M.MRAM[18][4] ),
    .I1(\mod.Data_Mem.F_M.MRAM[19][4] ),
    .S(_2301_),
    .Z(_2556_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _5936_ (.A1(_2366_),
    .A2(_2556_),
    .B(_2100_),
    .C(_2449_),
    .ZN(_2557_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5937_ (.I(_2402_),
    .Z(_2558_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5938_ (.I0(\mod.Data_Mem.F_M.MRAM[16][4] ),
    .I1(\mod.Data_Mem.F_M.MRAM[17][4] ),
    .S(_2189_),
    .Z(_2559_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5939_ (.I(_2396_),
    .Z(_2560_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5940_ (.A1(_2326_),
    .A2(\mod.Data_Mem.F_M.MRAM[21][4] ),
    .ZN(_2561_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5941_ (.A1(_2256_),
    .A2(\mod.Data_Mem.F_M.MRAM[20][4] ),
    .ZN(_2562_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _5942_ (.A1(_2560_),
    .A2(_2561_),
    .A3(_2562_),
    .ZN(_2563_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5943_ (.A1(_2558_),
    .A2(_2559_),
    .B(_2563_),
    .ZN(_2564_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5944_ (.I(_2065_),
    .Z(_2565_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _5945_ (.A1(_1533_),
    .A2(_2137_),
    .B1(_2557_),
    .B2(_2564_),
    .C(_2565_),
    .ZN(_2566_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5946_ (.I(_2283_),
    .Z(_2567_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5947_ (.I(_2102_),
    .Z(_2568_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _5948_ (.A1(_1778_),
    .A2(\mod.Data_Mem.F_M.MRAM[3][4] ),
    .Z(_2569_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _5949_ (.A1(_2567_),
    .A2(\mod.Data_Mem.F_M.MRAM[2][4] ),
    .B(_2568_),
    .C(_2569_),
    .ZN(_2570_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _5950_ (.A1(_2266_),
    .A2(\mod.Data_Mem.F_M.MRAM[4][4] ),
    .Z(_2571_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5951_ (.I(_2162_),
    .Z(_2572_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _5952_ (.A1(_2062_),
    .A2(\mod.Data_Mem.F_M.MRAM[5][4] ),
    .B(_2571_),
    .C(_2572_),
    .ZN(_2573_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _5953_ (.A1(_2266_),
    .A2(\mod.Data_Mem.F_M.MRAM[14][4] ),
    .Z(_2574_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _5954_ (.A1(_2506_),
    .A2(_1870_),
    .B(_2075_),
    .C(_2574_),
    .ZN(_2575_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _5955_ (.A1(_2410_),
    .A2(_2570_),
    .A3(_2573_),
    .A4(_2575_),
    .ZN(_2576_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _5956_ (.A1(_2531_),
    .A2(_2566_),
    .A3(_2576_),
    .ZN(_2577_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5957_ (.A1(_2534_),
    .A2(_2555_),
    .B1(_2577_),
    .B2(_2414_),
    .ZN(_0060_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5958_ (.I0(\mod.Data_Mem.F_M.MRAM[18][5] ),
    .I1(\mod.Data_Mem.F_M.MRAM[19][5] ),
    .S(_2161_),
    .Z(_2578_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _5959_ (.A1(_2457_),
    .A2(_2578_),
    .B(_1536_),
    .C(_2362_),
    .ZN(_2579_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5960_ (.I0(\mod.Data_Mem.F_M.MRAM[16][5] ),
    .I1(\mod.Data_Mem.F_M.MRAM[17][5] ),
    .S(_2283_),
    .Z(_2580_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5961_ (.A1(_2475_),
    .A2(\mod.Data_Mem.F_M.MRAM[21][5] ),
    .ZN(_2581_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5962_ (.A1(_2264_),
    .A2(\mod.Data_Mem.F_M.MRAM[20][5] ),
    .ZN(_2582_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _5963_ (.A1(_2397_),
    .A2(_2581_),
    .A3(_2582_),
    .ZN(_2583_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5964_ (.A1(_2558_),
    .A2(_2580_),
    .B(_2583_),
    .ZN(_2584_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _5965_ (.A1(_1627_),
    .A2(_2143_),
    .A3(_2145_),
    .ZN(_2585_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _5966_ (.A1(_2579_),
    .A2(_2584_),
    .B(_2585_),
    .C(_2263_),
    .ZN(_2586_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5967_ (.I(_2214_),
    .Z(_2587_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5968_ (.I(_1685_),
    .Z(_2588_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _5969_ (.A1(_2588_),
    .A2(\mod.Data_Mem.F_M.MRAM[4][5] ),
    .Z(_2589_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _5970_ (.A1(_2587_),
    .A2(\mod.Data_Mem.F_M.MRAM[5][5] ),
    .B(_2589_),
    .C(_2572_),
    .ZN(_2590_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5971_ (.I0(\mod.Data_Mem.F_M.MRAM[2][5] ),
    .I1(\mod.Data_Mem.F_M.MRAM[3][5] ),
    .S(_2540_),
    .Z(_2591_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5972_ (.I0(\mod.Data_Mem.F_M.MRAM[14][5] ),
    .I1(\mod.Data_Mem.F_M.MRAM[15][5] ),
    .S(_2528_),
    .Z(_2592_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5973_ (.A1(_2510_),
    .A2(_2591_),
    .B1(_2592_),
    .B2(_2565_),
    .ZN(_2593_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _5974_ (.A1(_2410_),
    .A2(_2590_),
    .A3(_2593_),
    .ZN(_2594_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _5975_ (.A1(_2531_),
    .A2(_2586_),
    .A3(_2594_),
    .ZN(_2595_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5976_ (.I(_2381_),
    .Z(_2596_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _5977_ (.A1(_1933_),
    .A2(\mod.Data_Mem.F_M.MRAM[783][5] ),
    .Z(_2597_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5978_ (.A1(_2385_),
    .A2(\mod.Data_Mem.F_M.MRAM[782][5] ),
    .B(_2597_),
    .ZN(_2598_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _5979_ (.A1(_2301_),
    .A2(\mod.Data_Mem.F_M.MRAM[773][5] ),
    .Z(_2599_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5980_ (.A1(_2343_),
    .A2(\mod.Data_Mem.F_M.MRAM[772][5] ),
    .B(_2599_),
    .ZN(_2600_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5981_ (.A1(_2596_),
    .A2(_2598_),
    .B1(_2600_),
    .B2(_2397_),
    .ZN(_2601_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5982_ (.I0(\mod.Data_Mem.F_M.MRAM[770][5] ),
    .I1(\mod.Data_Mem.F_M.MRAM[771][5] ),
    .S(_2522_),
    .Z(_2602_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5983_ (.A1(_2398_),
    .A2(_1934_),
    .ZN(_2603_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5984_ (.A1(_2424_),
    .A2(\mod.Data_Mem.F_M.MRAM[789][5] ),
    .B(_2603_),
    .ZN(_2604_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5985_ (.I0(\mod.Data_Mem.F_M.MRAM[786][5] ),
    .I1(\mod.Data_Mem.F_M.MRAM[787][5] ),
    .S(_1515_),
    .Z(_2605_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5986_ (.I0(\mod.Data_Mem.F_M.MRAM[784][5] ),
    .I1(\mod.Data_Mem.F_M.MRAM[785][5] ),
    .S(_1686_),
    .Z(_2606_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _5987_ (.A1(_2406_),
    .A2(_2605_),
    .B1(_2606_),
    .B2(_2403_),
    .ZN(_2607_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _5988_ (.A1(_2394_),
    .A2(_2142_),
    .B1(_2397_),
    .B2(_2604_),
    .C(_2607_),
    .ZN(_2608_));
 gf180mcu_fd_sc_mcu7t5v0__oai222_1 _5989_ (.A1(_1620_),
    .A2(_2601_),
    .B1(_2602_),
    .B2(_2104_),
    .C1(_2378_),
    .C2(_2608_),
    .ZN(_2609_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _5990_ (.A1(_2079_),
    .A2(_2609_),
    .Z(_2610_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5991_ (.A1(_2414_),
    .A2(_2595_),
    .B(_2610_),
    .ZN(_0061_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5992_ (.I(_2560_),
    .Z(_2611_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _5993_ (.A1(_2588_),
    .A2(\mod.Data_Mem.F_M.MRAM[789][6] ),
    .Z(_2612_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5994_ (.A1(_2587_),
    .A2(\mod.Data_Mem.F_M.MRAM[788][6] ),
    .B(_2612_),
    .ZN(_2613_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5995_ (.A1(_2214_),
    .A2(\mod.Data_Mem.F_M.MRAM[786][6] ),
    .ZN(_2614_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5996_ (.A1(_2313_),
    .A2(_2013_),
    .B(_2614_),
    .ZN(_2615_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5997_ (.I0(\mod.Data_Mem.F_M.MRAM[784][6] ),
    .I1(\mod.Data_Mem.F_M.MRAM[785][6] ),
    .S(_2331_),
    .Z(_2616_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _5998_ (.A1(_2464_),
    .A2(_2615_),
    .B1(_2616_),
    .B2(_2539_),
    .ZN(_2617_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _5999_ (.A1(_2535_),
    .A2(_2150_),
    .B1(_2611_),
    .B2(_2613_),
    .C(_2617_),
    .ZN(_2618_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6000_ (.I(_1778_),
    .Z(_2619_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6001_ (.I(_1681_),
    .Z(_2620_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _6002_ (.A1(_2620_),
    .A2(\mod.Data_Mem.F_M.MRAM[783][6] ),
    .Z(_2621_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6003_ (.A1(_2619_),
    .A2(\mod.Data_Mem.F_M.MRAM[782][6] ),
    .B(_2621_),
    .ZN(_2622_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _6004_ (.A1(_2588_),
    .A2(\mod.Data_Mem.F_M.MRAM[773][6] ),
    .Z(_2623_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6005_ (.A1(_2062_),
    .A2(\mod.Data_Mem.F_M.MRAM[772][6] ),
    .B(_2623_),
    .ZN(_2624_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6006_ (.A1(_2535_),
    .A2(_2622_),
    .B1(_2624_),
    .B2(_2611_),
    .ZN(_2625_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6007_ (.I(_1757_),
    .Z(_2626_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6008_ (.I0(\mod.Data_Mem.F_M.MRAM[770][6] ),
    .I1(\mod.Data_Mem.F_M.MRAM[771][6] ),
    .S(_2275_),
    .Z(_2627_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6009_ (.A1(_2104_),
    .A2(_2627_),
    .ZN(_2628_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6010_ (.A1(_2413_),
    .A2(_2628_),
    .ZN(_2629_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _6011_ (.A1(_2379_),
    .A2(_2618_),
    .B1(_2625_),
    .B2(_2626_),
    .C(_2629_),
    .ZN(_2630_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6012_ (.I0(\mod.Data_Mem.F_M.MRAM[16][6] ),
    .I1(\mod.Data_Mem.F_M.MRAM[17][6] ),
    .S(_2418_),
    .Z(_2631_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6013_ (.A1(_2549_),
    .A2(\mod.Data_Mem.F_M.MRAM[20][6] ),
    .ZN(_2632_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6014_ (.A1(_2512_),
    .A2(\mod.Data_Mem.F_M.MRAM[21][6] ),
    .ZN(_2633_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6015_ (.A1(_2548_),
    .A2(_2632_),
    .A3(_2633_),
    .ZN(_2634_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _6016_ (.A1(_1685_),
    .A2(\mod.Data_Mem.F_M.MRAM[19][6] ),
    .Z(_2635_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6017_ (.A1(_2061_),
    .A2(\mod.Data_Mem.F_M.MRAM[18][6] ),
    .B(_2635_),
    .ZN(_2636_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6018_ (.A1(_2352_),
    .A2(_2636_),
    .B(_2354_),
    .ZN(_2637_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _6019_ (.A1(_2558_),
    .A2(_2631_),
    .B(_2634_),
    .C(_2637_),
    .ZN(_2638_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _6020_ (.A1(_2185_),
    .A2(_2148_),
    .B(_2638_),
    .C(_2263_),
    .ZN(_2639_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _6021_ (.A1(_2345_),
    .A2(\mod.Data_Mem.F_M.MRAM[4][6] ),
    .Z(_2640_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _6022_ (.A1(_2587_),
    .A2(\mod.Data_Mem.F_M.MRAM[5][6] ),
    .B(_2640_),
    .C(_2091_),
    .ZN(_2641_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6023_ (.I(_2388_),
    .Z(_2642_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6024_ (.I0(\mod.Data_Mem.F_M.MRAM[2][6] ),
    .I1(\mod.Data_Mem.F_M.MRAM[3][6] ),
    .S(_2528_),
    .Z(_2643_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6025_ (.I0(\mod.Data_Mem.F_M.MRAM[14][6] ),
    .I1(\mod.Data_Mem.F_M.MRAM[15][6] ),
    .S(_2360_),
    .Z(_2644_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6026_ (.A1(_2642_),
    .A2(_2643_),
    .B1(_2644_),
    .B2(_2565_),
    .ZN(_2645_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6027_ (.A1(_2416_),
    .A2(_2641_),
    .A3(_2645_),
    .ZN(_2646_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _6028_ (.A1(_1670_),
    .A2(_2118_),
    .A3(_2639_),
    .A4(_2646_),
    .ZN(_2647_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6029_ (.A1(_2630_),
    .A2(_2647_),
    .ZN(_0062_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _6030_ (.A1(_2428_),
    .A2(\mod.Data_Mem.F_M.MRAM[789][7] ),
    .Z(_2648_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6031_ (.A1(_2506_),
    .A2(\mod.Data_Mem.F_M.MRAM[788][7] ),
    .B(_2648_),
    .ZN(_2649_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6032_ (.I0(\mod.Data_Mem.F_M.MRAM[784][7] ),
    .I1(\mod.Data_Mem.F_M.MRAM[785][7] ),
    .S(_2331_),
    .Z(_2650_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6033_ (.A1(_2097_),
    .A2(\mod.Data_Mem.F_M.MRAM[786][7] ),
    .ZN(_2651_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6034_ (.A1(_2549_),
    .A2(_2049_),
    .B(_2651_),
    .ZN(_2652_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _6035_ (.A1(_2539_),
    .A2(_2650_),
    .B1(_2652_),
    .B2(_2435_),
    .ZN(_2653_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _6036_ (.A1(_2535_),
    .A2(_2156_),
    .B1(_2536_),
    .B2(_2649_),
    .C(_2653_),
    .ZN(_2654_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6037_ (.I0(\mod.Data_Mem.F_M.MRAM[782][7] ),
    .I1(\mod.Data_Mem.F_M.MRAM[783][7] ),
    .S(_2326_),
    .Z(_2655_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6038_ (.I0(\mod.Data_Mem.F_M.MRAM[770][7] ),
    .I1(\mod.Data_Mem.F_M.MRAM[771][7] ),
    .S(_2339_),
    .Z(_2656_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6039_ (.A1(_2288_),
    .A2(\mod.Data_Mem.F_M.MRAM[773][7] ),
    .ZN(_2657_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6040_ (.A1(_2549_),
    .A2(\mod.Data_Mem.F_M.MRAM[772][7] ),
    .ZN(_2658_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6041_ (.A1(_2548_),
    .A2(_2657_),
    .A3(_2658_),
    .ZN(_2659_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _6042_ (.A1(_2423_),
    .A2(_2655_),
    .B1(_2656_),
    .B2(_2464_),
    .C(_2659_),
    .ZN(_2660_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6043_ (.A1(_2434_),
    .A2(_2660_),
    .ZN(_2661_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6044_ (.A1(_2379_),
    .A2(_2654_),
    .B(_2661_),
    .ZN(_2662_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6045_ (.I0(\mod.Data_Mem.F_M.MRAM[16][7] ),
    .I1(\mod.Data_Mem.F_M.MRAM[17][7] ),
    .S(_2540_),
    .Z(_2663_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6046_ (.A1(_2620_),
    .A2(\mod.Data_Mem.F_M.MRAM[21][7] ),
    .ZN(_2664_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6047_ (.A1(_2214_),
    .A2(\mod.Data_Mem.F_M.MRAM[20][7] ),
    .ZN(_2665_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6048_ (.A1(_2560_),
    .A2(_2664_),
    .A3(_2665_),
    .ZN(_2666_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _6049_ (.A1(_1612_),
    .A2(\mod.Data_Mem.F_M.MRAM[19][7] ),
    .Z(_2667_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6050_ (.A1(_2129_),
    .A2(\mod.Data_Mem.F_M.MRAM[18][7] ),
    .B(_2667_),
    .ZN(_2668_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6051_ (.A1(_2352_),
    .A2(_2668_),
    .B(_2354_),
    .ZN(_2669_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _6052_ (.A1(_2539_),
    .A2(_2663_),
    .B(_2666_),
    .C(_2669_),
    .ZN(_2670_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _6053_ (.A1(_2185_),
    .A2(_2154_),
    .B(_2670_),
    .C(_2263_),
    .ZN(_2671_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6054_ (.I(_2495_),
    .Z(_2672_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6055_ (.I0(\mod.Data_Mem.F_M.MRAM[2][7] ),
    .I1(\mod.Data_Mem.F_M.MRAM[3][7] ),
    .S(_1769_),
    .Z(_2673_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6056_ (.A1(_2672_),
    .A2(_2673_),
    .ZN(_2674_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _6057_ (.A1(_2288_),
    .A2(\mod.Data_Mem.F_M.MRAM[4][7] ),
    .Z(_2675_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _6058_ (.A1(_2062_),
    .A2(\mod.Data_Mem.F_M.MRAM[5][7] ),
    .B(_2675_),
    .C(_2572_),
    .ZN(_2676_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6059_ (.I0(\mod.Data_Mem.F_M.MRAM[14][7] ),
    .I1(\mod.Data_Mem.F_M.MRAM[15][7] ),
    .S(_2295_),
    .Z(_2677_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6060_ (.A1(_2565_),
    .A2(_2677_),
    .ZN(_2678_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _6061_ (.A1(_2410_),
    .A2(_2674_),
    .A3(_2676_),
    .A4(_2678_),
    .ZN(_2679_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6062_ (.A1(_2531_),
    .A2(_2671_),
    .A3(_2679_),
    .ZN(_2680_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6063_ (.A1(_2534_),
    .A2(_2662_),
    .B1(_2680_),
    .B2(_2414_),
    .ZN(_0063_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _6064_ (.A1(_1840_),
    .A2(_2402_),
    .B(_1535_),
    .ZN(_2681_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6065_ (.I(_2681_),
    .Z(_2682_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _6066_ (.A1(_2517_),
    .A2(\mod.Data_Mem.F_M.MRAM[782][0] ),
    .B1(\mod.Data_Mem.F_M.MRAM[783][0] ),
    .B2(_2567_),
    .ZN(_2683_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6067_ (.A1(_2682_),
    .A2(_2683_),
    .ZN(_2684_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _6068_ (.A1(_1676_),
    .A2(_2375_),
    .B(_1495_),
    .ZN(_2685_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6069_ (.I(_2685_),
    .Z(_2686_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6070_ (.I(_2686_),
    .Z(_2687_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6071_ (.A1(_2172_),
    .A2(_2687_),
    .B(_1729_),
    .ZN(_2688_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6072_ (.I(_2681_),
    .Z(_2689_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6073_ (.A1(\mod.Data_Mem.F_M.MRAM[797][0] ),
    .A2(_2689_),
    .ZN(_2690_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6074_ (.I(_2685_),
    .Z(_2691_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6075_ (.I(_2691_),
    .Z(_2692_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6076_ (.A1(\mod.Data_Mem.F_M.MRAM[781][0] ),
    .A2(_2692_),
    .ZN(_2693_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6077_ (.A1(_2087_),
    .A2(_2690_),
    .A3(_2693_),
    .ZN(_2694_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _6078_ (.A1(_2684_),
    .A2(_2688_),
    .B(_1726_),
    .C(_2694_),
    .ZN(_2695_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6079_ (.I(_2295_),
    .Z(_2696_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6080_ (.A1(_2696_),
    .A2(\mod.Data_Mem.F_M.MRAM[14][0] ),
    .B1(\mod.Data_Mem.F_M.MRAM[15][0] ),
    .B2(_2517_),
    .ZN(_2697_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6081_ (.I(_1756_),
    .Z(_2698_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _6082_ (.A1(\mod.Data_Mem.F_M.MRAM[13][0] ),
    .A2(_2087_),
    .B1(_2212_),
    .B2(\mod.Data_Mem.F_M.MRAM[12][0] ),
    .C(_2698_),
    .ZN(_2699_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6083_ (.A1(_1802_),
    .A2(_2697_),
    .B(_2699_),
    .ZN(_2700_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _6084_ (.A1(_2081_),
    .A2(_1497_),
    .B1(_2165_),
    .B2(_1620_),
    .C(_1965_),
    .ZN(_2701_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6085_ (.A1(_2209_),
    .A2(_2201_),
    .ZN(_2702_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6086_ (.I(_2702_),
    .Z(_2703_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6087_ (.A1(_2700_),
    .A2(_2701_),
    .B(_2703_),
    .ZN(_2704_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6088_ (.A1(_2012_),
    .A2(_1610_),
    .ZN(_2705_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6089_ (.A1(_1494_),
    .A2(_1542_),
    .Z(_2706_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6090_ (.I(_2706_),
    .Z(_2707_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6091_ (.I(_2707_),
    .Z(_2708_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6092_ (.A1(_1764_),
    .A2(_1613_),
    .ZN(_2709_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6093_ (.A1(_2705_),
    .A2(_2708_),
    .A3(_2709_),
    .ZN(_2710_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6094_ (.A1(_2326_),
    .A2(\mod.Data_Mem.F_M.MRAM[790][0] ),
    .B1(\mod.Data_Mem.F_M.MRAM[791][0] ),
    .B2(_2116_),
    .ZN(_2711_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6095_ (.A1(_2196_),
    .A2(_1604_),
    .ZN(_2712_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6096_ (.A1(_1500_),
    .A2(_1541_),
    .Z(_2713_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6097_ (.I(_2713_),
    .Z(_2714_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6098_ (.I(_2714_),
    .Z(_2715_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _6099_ (.A1(_2195_),
    .A2(_2711_),
    .B(_2712_),
    .C(_2715_),
    .ZN(_2716_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6100_ (.A1(_2710_),
    .A2(_2689_),
    .A3(_2716_),
    .ZN(_2717_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6101_ (.I(_2707_),
    .Z(_2718_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6102_ (.A1(_2186_),
    .A2(_1582_),
    .ZN(_2719_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6103_ (.A1(_1764_),
    .A2(_1589_),
    .ZN(_2720_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6104_ (.A1(_2718_),
    .A2(_2719_),
    .A3(_2720_),
    .ZN(_2721_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6105_ (.A1(_2620_),
    .A2(\mod.Data_Mem.F_M.MRAM[774][0] ),
    .B1(\mod.Data_Mem.F_M.MRAM[775][0] ),
    .B2(_2162_),
    .ZN(_2722_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6106_ (.I(_1737_),
    .Z(_2723_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6107_ (.A1(_2723_),
    .A2(_1569_),
    .ZN(_2724_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _6108_ (.A1(_1640_),
    .A2(_2722_),
    .B(_2724_),
    .C(_2715_),
    .ZN(_2725_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6109_ (.A1(_2692_),
    .A2(_2721_),
    .A3(_2725_),
    .ZN(_2726_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6110_ (.A1(_2185_),
    .A2(_2717_),
    .A3(_2726_),
    .ZN(_2727_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6111_ (.I(_1691_),
    .Z(_2728_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _6112_ (.A1(_2540_),
    .A2(\mod.Data_Mem.F_M.MRAM[2][0] ),
    .Z(_2729_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _6113_ (.A1(_2728_),
    .A2(\mod.Data_Mem.F_M.MRAM[3][0] ),
    .B(_1805_),
    .C(_2729_),
    .ZN(_2730_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _6114_ (.A1(\mod.Data_Mem.F_M.MRAM[1][0] ),
    .A2(_1539_),
    .B1(_1809_),
    .B2(\mod.Data_Mem.F_M.MRAM[0][0] ),
    .C(_2708_),
    .ZN(_2731_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6115_ (.I0(\mod.Data_Mem.F_M.MRAM[7][0] ),
    .I1(\mod.Data_Mem.F_M.MRAM[6][0] ),
    .S(_1707_),
    .Z(_2732_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6116_ (.I(_2714_),
    .Z(_2733_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _6117_ (.A1(_1540_),
    .A2(_1505_),
    .B1(_1575_),
    .B2(_2732_),
    .C(_2733_),
    .ZN(_2734_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _6118_ (.A1(_2373_),
    .A2(_2687_),
    .B1(_2730_),
    .B2(_2731_),
    .C(_2734_),
    .ZN(_2735_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6119_ (.I0(\mod.Data_Mem.F_M.MRAM[23][0] ),
    .I1(\mod.Data_Mem.F_M.MRAM[22][0] ),
    .S(_1782_),
    .Z(_2736_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _6120_ (.A1(_1505_),
    .A2(_1511_),
    .B1(_2736_),
    .B2(_1575_),
    .C(_2733_),
    .ZN(_2737_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6121_ (.A1(_2373_),
    .A2(_2691_),
    .ZN(_2738_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6122_ (.I(_2706_),
    .Z(_2739_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _6123_ (.A1(_1795_),
    .A2(_1516_),
    .B1(_1520_),
    .B2(_1713_),
    .C(_2739_),
    .ZN(_2740_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _6124_ (.A1(_2738_),
    .A2(_2740_),
    .Z(_2741_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _6125_ (.A1(_2696_),
    .A2(_1497_),
    .B1(_2737_),
    .B2(_2741_),
    .C(_1625_),
    .ZN(_2742_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _6126_ (.A1(_2366_),
    .A2(_2195_),
    .ZN(_2743_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _6127_ (.A1(_1726_),
    .A2(_2727_),
    .B1(_2735_),
    .B2(_2742_),
    .C(_2743_),
    .ZN(_2744_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6128_ (.A1(_2695_),
    .A2(_2704_),
    .B(_2744_),
    .ZN(_0064_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6129_ (.A1(_2619_),
    .A2(\mod.Data_Mem.F_M.MRAM[783][1] ),
    .B1(\mod.Data_Mem.F_M.MRAM[782][1] ),
    .B2(_2089_),
    .ZN(_2745_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _6130_ (.A1(\mod.Data_Mem.F_M.MRAM[781][1] ),
    .A2(_2200_),
    .B1(_1809_),
    .B2(\mod.Data_Mem.F_M.MRAM[780][1] ),
    .ZN(_2746_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6131_ (.A1(_2169_),
    .A2(_2745_),
    .B(_2746_),
    .ZN(_2747_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6132_ (.A1(_2183_),
    .A2(_2689_),
    .ZN(_2748_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _6133_ (.A1(_2682_),
    .A2(_2747_),
    .B(_2748_),
    .C(_2084_),
    .ZN(_2749_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6134_ (.I(_2685_),
    .Z(_2750_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6135_ (.I(_1538_),
    .Z(_2751_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6136_ (.I(_1564_),
    .Z(_2752_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _6137_ (.A1(_2009_),
    .A2(\mod.Data_Mem.F_M.MRAM[14][1] ),
    .B1(\mod.Data_Mem.F_M.MRAM[15][1] ),
    .B2(_1968_),
    .ZN(_2753_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6138_ (.A1(_2752_),
    .A2(_2753_),
    .ZN(_2754_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _6139_ (.A1(\mod.Data_Mem.F_M.MRAM[13][1] ),
    .A2(_2751_),
    .B1(_2157_),
    .B2(\mod.Data_Mem.F_M.MRAM[12][1] ),
    .C(_2754_),
    .ZN(_2755_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _6140_ (.A1(_2750_),
    .A2(_2755_),
    .Z(_2756_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _6141_ (.A1(_2192_),
    .A2(_2689_),
    .B(_2756_),
    .C(_1625_),
    .ZN(_2757_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6142_ (.A1(_2703_),
    .A2(_2757_),
    .ZN(_2758_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6143_ (.I(_2691_),
    .Z(_2759_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6144_ (.A1(_2360_),
    .A2(\mod.Data_Mem.F_M.MRAM[6][1] ),
    .B1(\mod.Data_Mem.F_M.MRAM[7][1] ),
    .B2(_2188_),
    .ZN(_2760_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6145_ (.I(_1573_),
    .Z(_2761_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6146_ (.A1(_2761_),
    .A2(_1637_),
    .ZN(_2762_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6147_ (.I(_2713_),
    .Z(_2763_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _6148_ (.A1(_1640_),
    .A2(_2760_),
    .B(_2762_),
    .C(_2763_),
    .ZN(_2764_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6149_ (.I(_2706_),
    .Z(_2765_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6150_ (.A1(_1742_),
    .A2(_1648_),
    .ZN(_2766_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6151_ (.A1(_2180_),
    .A2(_1649_),
    .ZN(_2767_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6152_ (.A1(_2765_),
    .A2(_2766_),
    .A3(_2767_),
    .ZN(_2768_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6153_ (.A1(_2759_),
    .A2(_2764_),
    .A3(_2768_),
    .ZN(_2769_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6154_ (.A1(_1751_),
    .A2(_1659_),
    .ZN(_2770_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6155_ (.A1(_1910_),
    .A2(_1656_),
    .ZN(_2771_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6156_ (.A1(_2765_),
    .A2(_2770_),
    .A3(_2771_),
    .ZN(_2772_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6157_ (.A1(_2425_),
    .A2(\mod.Data_Mem.F_M.MRAM[22][1] ),
    .B1(\mod.Data_Mem.F_M.MRAM[23][1] ),
    .B2(_2188_),
    .ZN(_2773_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6158_ (.A1(_2761_),
    .A2(_1665_),
    .ZN(_2774_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6159_ (.I(_2713_),
    .Z(_2775_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _6160_ (.A1(_1661_),
    .A2(_2773_),
    .B(_2774_),
    .C(_2775_),
    .ZN(_2776_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6161_ (.A1(_2681_),
    .A2(_2772_),
    .A3(_2776_),
    .ZN(_2777_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6162_ (.A1(_2769_),
    .A2(_2777_),
    .ZN(_2778_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6163_ (.I(_2707_),
    .Z(_2779_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6164_ (.A1(_1555_),
    .A2(_1702_),
    .B1(_1703_),
    .B2(_1566_),
    .ZN(_2780_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6165_ (.A1(_1706_),
    .A2(_1718_),
    .ZN(_2781_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6166_ (.A1(_1730_),
    .A2(_1711_),
    .ZN(_2782_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6167_ (.A1(_2708_),
    .A2(_2781_),
    .A3(_2782_),
    .ZN(_2783_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _6168_ (.A1(_2779_),
    .A2(_2780_),
    .B(_2783_),
    .C(_2692_),
    .ZN(_2784_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6169_ (.A1(_2186_),
    .A2(_1694_),
    .ZN(_2785_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6170_ (.A1(_2196_),
    .A2(_1689_),
    .B(_2739_),
    .ZN(_2786_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6171_ (.A1(_1645_),
    .A2(_1680_),
    .ZN(_2787_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6172_ (.A1(_1734_),
    .A2(_1684_),
    .B(_2775_),
    .ZN(_2788_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _6173_ (.A1(_2785_),
    .A2(_2786_),
    .B1(_2787_),
    .B2(_2788_),
    .C(_2750_),
    .ZN(_2789_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6174_ (.A1(_1898_),
    .A2(_2789_),
    .ZN(_2790_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _6175_ (.A1(_1670_),
    .A2(_2778_),
    .B1(_2784_),
    .B2(_2790_),
    .C(_2743_),
    .ZN(_2791_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _6176_ (.A1(_2749_),
    .A2(_2758_),
    .B(_2791_),
    .C(_2374_),
    .ZN(_0065_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6177_ (.A1(_2199_),
    .A2(_2682_),
    .ZN(_2792_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6178_ (.A1(_2319_),
    .A2(\mod.Data_Mem.F_M.MRAM[783][2] ),
    .B1(\mod.Data_Mem.F_M.MRAM[782][2] ),
    .B2(_2311_),
    .ZN(_2793_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6179_ (.A1(_1585_),
    .A2(_2793_),
    .ZN(_2794_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _6180_ (.A1(\mod.Data_Mem.F_M.MRAM[781][2] ),
    .A2(_2200_),
    .B1(_2202_),
    .B2(\mod.Data_Mem.F_M.MRAM[780][2] ),
    .C(_2794_),
    .ZN(_2795_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6181_ (.A1(_2687_),
    .A2(_2795_),
    .ZN(_2796_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6182_ (.A1(_2073_),
    .A2(_2792_),
    .A3(_2796_),
    .ZN(_2797_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6183_ (.A1(_2206_),
    .A2(_2682_),
    .ZN(_2798_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6184_ (.A1(_2070_),
    .A2(\mod.Data_Mem.F_M.MRAM[14][2] ),
    .B1(\mod.Data_Mem.F_M.MRAM[15][2] ),
    .B2(_2203_),
    .ZN(_2799_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6185_ (.A1(_1834_),
    .A2(_2799_),
    .ZN(_2800_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _6186_ (.A1(\mod.Data_Mem.F_M.MRAM[13][2] ),
    .A2(_2200_),
    .B1(_2202_),
    .B2(\mod.Data_Mem.F_M.MRAM[12][2] ),
    .C(_2800_),
    .ZN(_2801_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6187_ (.A1(_2687_),
    .A2(_2801_),
    .B(_1965_),
    .ZN(_2802_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6188_ (.A1(_2798_),
    .A2(_2802_),
    .B(_2703_),
    .ZN(_2803_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6189_ (.A1(_2360_),
    .A2(\mod.Data_Mem.F_M.MRAM[6][2] ),
    .B1(\mod.Data_Mem.F_M.MRAM[7][2] ),
    .B2(_2188_),
    .ZN(_2804_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6190_ (.A1(_2761_),
    .A2(_1731_),
    .ZN(_2805_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _6191_ (.A1(_1661_),
    .A2(_2804_),
    .B(_2805_),
    .C(_2763_),
    .ZN(_2806_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6192_ (.A1(_1742_),
    .A2(_1739_),
    .ZN(_2807_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6193_ (.A1(_2180_),
    .A2(_1735_),
    .ZN(_2808_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6194_ (.A1(_2765_),
    .A2(_2807_),
    .A3(_2808_),
    .ZN(_2809_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6195_ (.A1(_2759_),
    .A2(_2806_),
    .A3(_2809_),
    .ZN(_2810_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6196_ (.A1(_1751_),
    .A2(_1747_),
    .ZN(_2811_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6197_ (.A1(_1910_),
    .A2(_1743_),
    .ZN(_2812_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6198_ (.A1(_2765_),
    .A2(_2811_),
    .A3(_2812_),
    .ZN(_2813_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6199_ (.A1(_2425_),
    .A2(\mod.Data_Mem.F_M.MRAM[22][2] ),
    .B1(\mod.Data_Mem.F_M.MRAM[23][2] ),
    .B2(_2448_),
    .ZN(_2814_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6200_ (.A1(_2761_),
    .A2(_1752_),
    .ZN(_2815_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _6201_ (.A1(_1661_),
    .A2(_2814_),
    .B(_2815_),
    .C(_2775_),
    .ZN(_2816_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6202_ (.A1(_2681_),
    .A2(_2813_),
    .A3(_2816_),
    .ZN(_2817_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6203_ (.A1(_2810_),
    .A2(_2817_),
    .ZN(_2818_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6204_ (.A1(_1566_),
    .A2(_1761_),
    .B1(_1762_),
    .B2(_1555_),
    .ZN(_2819_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6205_ (.A1(_1706_),
    .A2(_1772_),
    .ZN(_2820_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6206_ (.A1(_1730_),
    .A2(_1767_),
    .ZN(_2821_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6207_ (.A1(_2708_),
    .A2(_2820_),
    .A3(_2821_),
    .ZN(_2822_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _6208_ (.A1(_2779_),
    .A2(_2819_),
    .B(_2822_),
    .C(_2692_),
    .ZN(_2823_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6209_ (.A1(_2186_),
    .A2(_1781_),
    .ZN(_2824_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6210_ (.A1(_2196_),
    .A2(_1786_),
    .B(_2739_),
    .ZN(_2825_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6211_ (.A1(_1706_),
    .A2(_1794_),
    .ZN(_2826_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6212_ (.A1(_1734_),
    .A2(_1789_),
    .B(_2775_),
    .ZN(_2827_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _6213_ (.A1(_2824_),
    .A2(_2825_),
    .B1(_2826_),
    .B2(_2827_),
    .C(_2686_),
    .ZN(_2828_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6214_ (.A1(_1898_),
    .A2(_2828_),
    .ZN(_2829_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _6215_ (.A1(_1800_),
    .A2(_2818_),
    .B1(_2823_),
    .B2(_2829_),
    .C(_2743_),
    .ZN(_2830_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _6216_ (.A1(_2797_),
    .A2(_2803_),
    .B(_2830_),
    .C(_2374_),
    .ZN(_0066_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6217_ (.I(_2107_),
    .Z(_2831_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6218_ (.A1(_2212_),
    .A2(_2219_),
    .B(_2508_),
    .ZN(_2832_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6219_ (.A1(_2567_),
    .A2(_2572_),
    .A3(\mod.Data_Mem.F_M.MRAM[20][3] ),
    .ZN(_2833_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6220_ (.A1(_2832_),
    .A2(_2833_),
    .ZN(_2834_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _6221_ (.I0(\mod.Data_Mem.F_M.MRAM[1][3] ),
    .I1(\mod.Data_Mem.F_M.MRAM[2][3] ),
    .I2(\mod.Data_Mem.F_M.MRAM[3][3] ),
    .I3(\mod.Data_Mem.F_M.MRAM[4][3] ),
    .S0(_2588_),
    .S1(_2449_),
    .Z(_2835_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _6222_ (.A1(_1734_),
    .A2(_1819_),
    .Z(_2836_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6223_ (.A1(_2714_),
    .A2(_2685_),
    .ZN(_2837_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _6224_ (.A1(_1931_),
    .A2(_1817_),
    .B(_2836_),
    .C(_2837_),
    .ZN(_2838_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6225_ (.A1(_2217_),
    .A2(\mod.Data_Mem.F_M.MRAM[14][3] ),
    .B1(\mod.Data_Mem.F_M.MRAM[15][3] ),
    .B2(_2319_),
    .ZN(_2839_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6226_ (.A1(_1585_),
    .A2(_2839_),
    .ZN(_2840_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6227_ (.A1(_1619_),
    .A2(_2702_),
    .ZN(_2841_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _6228_ (.A1(\mod.Data_Mem.F_M.MRAM[13][3] ),
    .A2(_1729_),
    .B(_2840_),
    .C(_2841_),
    .ZN(_2842_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6229_ (.A1(_2838_),
    .A2(_2842_),
    .ZN(_2843_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _6230_ (.A1(_2831_),
    .A2(_2834_),
    .B1(_2835_),
    .B2(_2093_),
    .C(_2843_),
    .ZN(_2844_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6231_ (.A1(_2169_),
    .A2(_1837_),
    .ZN(_2845_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6232_ (.I(_2714_),
    .Z(_2846_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6233_ (.A1(_1802_),
    .A2(_1832_),
    .B(_2846_),
    .ZN(_2847_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _6234_ (.A1(_2723_),
    .A2(_1830_),
    .Z(_2848_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _6235_ (.A1(_2160_),
    .A2(_1827_),
    .B(_2718_),
    .C(_2848_),
    .ZN(_2849_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _6236_ (.A1(_2845_),
    .A2(_2847_),
    .B(_2738_),
    .C(_2849_),
    .ZN(_2850_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6237_ (.A1(_1931_),
    .A2(_1848_),
    .ZN(_2851_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6238_ (.A1(_2160_),
    .A2(_1842_),
    .ZN(_2852_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6239_ (.A1(_2846_),
    .A2(_2851_),
    .A3(_2852_),
    .ZN(_2853_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6240_ (.A1(_2160_),
    .A2(_1853_),
    .ZN(_2854_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6241_ (.A1(_1931_),
    .A2(_1857_),
    .B(_2733_),
    .ZN(_2855_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6242_ (.A1(_2854_),
    .A2(_2855_),
    .B(_2738_),
    .ZN(_2856_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6243_ (.A1(_2853_),
    .A2(_2856_),
    .B(_2743_),
    .ZN(_2857_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6244_ (.I(\mod.Data_Mem.F_M.MRAM[781][3] ),
    .ZN(_2858_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6245_ (.A1(_2129_),
    .A2(\mod.Data_Mem.F_M.MRAM[783][3] ),
    .B1(\mod.Data_Mem.F_M.MRAM[782][3] ),
    .B2(_2070_),
    .ZN(_2859_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6246_ (.A1(_2858_),
    .A2(_2221_),
    .B1(_1664_),
    .B2(_2859_),
    .ZN(_2860_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _6247_ (.A1(_2107_),
    .A2(_2860_),
    .B(_2202_),
    .C(_2210_),
    .ZN(_2861_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6248_ (.A1(_2108_),
    .A2(_2224_),
    .B(_2861_),
    .ZN(_2862_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6249_ (.A1(_2850_),
    .A2(_2857_),
    .B(_2862_),
    .ZN(_2863_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6250_ (.A1(_2212_),
    .A2(_1627_),
    .ZN(_2864_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6251_ (.A1(_2079_),
    .A2(_2864_),
    .ZN(_2865_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _6252_ (.A1(_2534_),
    .A2(_2844_),
    .B1(_2863_),
    .B2(_2865_),
    .ZN(_0067_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6253_ (.I(_2374_),
    .Z(_2866_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6254_ (.I(_2702_),
    .Z(_2867_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6255_ (.I(_2867_),
    .Z(_2868_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6256_ (.I(_2686_),
    .Z(_2869_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6257_ (.I(_1574_),
    .Z(_2870_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6258_ (.A1(_2870_),
    .A2(_1874_),
    .ZN(_2871_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6259_ (.I(_1663_),
    .Z(_2872_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6260_ (.I(_2706_),
    .Z(_2873_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6261_ (.A1(_2872_),
    .A2(_1876_),
    .B(_2873_),
    .ZN(_2874_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6262_ (.A1(_1655_),
    .A2(_1880_),
    .ZN(_2875_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6263_ (.I(_1737_),
    .Z(_2876_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6264_ (.A1(_2876_),
    .A2(_1878_),
    .B(_2715_),
    .ZN(_2877_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6265_ (.A1(_2871_),
    .A2(_2874_),
    .B1(_2875_),
    .B2(_2877_),
    .ZN(_2878_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6266_ (.A1(_2869_),
    .A2(_2878_),
    .ZN(_2879_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6267_ (.I0(_1889_),
    .I1(_1891_),
    .S(_2723_),
    .Z(_2880_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6268_ (.A1(_2707_),
    .A2(_2691_),
    .ZN(_2881_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6269_ (.I(_2881_),
    .Z(_2882_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6270_ (.I0(_1895_),
    .I1(_1893_),
    .S(_1742_),
    .Z(_2883_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6271_ (.I(_2837_),
    .Z(_2884_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _6272_ (.A1(_2880_),
    .A2(_2882_),
    .B1(_2883_),
    .B2(_2884_),
    .C(_1490_),
    .ZN(_2885_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6273_ (.I(_2686_),
    .Z(_2886_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6274_ (.A1(_1941_),
    .A2(_1904_),
    .ZN(_2887_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6275_ (.A1(_2872_),
    .A2(_1905_),
    .ZN(_2888_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6276_ (.A1(_2846_),
    .A2(_2887_),
    .A3(_2888_),
    .ZN(_2889_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6277_ (.A1(_1826_),
    .A2(_1909_),
    .ZN(_2890_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6278_ (.I(_2228_),
    .Z(_2891_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6279_ (.A1(_2891_),
    .A2(_1907_),
    .ZN(_2892_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6280_ (.A1(_2718_),
    .A2(_2890_),
    .A3(_2892_),
    .ZN(_2893_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6281_ (.A1(_2886_),
    .A2(_2889_),
    .A3(_2893_),
    .ZN(_2894_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6282_ (.I(_2881_),
    .Z(_2895_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _6283_ (.I0(\mod.Data_Mem.F_M.MRAM[789][4] ),
    .I1(\mod.Data_Mem.F_M.MRAM[791][4] ),
    .I2(\mod.Data_Mem.F_M.MRAM[790][4] ),
    .I3(\mod.Data_Mem.F_M.MRAM[788][4] ),
    .S0(_2448_),
    .S1(_2383_),
    .Z(_2896_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6284_ (.I0(_1921_),
    .I1(_1922_),
    .S(_2044_),
    .Z(_2897_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6285_ (.I(_2837_),
    .Z(_2898_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _6286_ (.A1(_2895_),
    .A2(_2896_),
    .B1(_2897_),
    .B2(_2898_),
    .C(_1866_),
    .ZN(_2899_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6287_ (.A1(_2879_),
    .A2(_2885_),
    .B1(_2894_),
    .B2(_2899_),
    .ZN(_2900_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6288_ (.I(_1537_),
    .Z(_2901_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6289_ (.I(_1543_),
    .Z(_2902_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6290_ (.I(_1564_),
    .Z(_2903_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6291_ (.I(_2059_),
    .Z(_2904_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6292_ (.I(_1493_),
    .Z(_2905_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6293_ (.A1(_2904_),
    .A2(\mod.Data_Mem.F_M.MRAM[15][4] ),
    .B1(\mod.Data_Mem.F_M.MRAM[14][4] ),
    .B2(_2905_),
    .ZN(_2906_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6294_ (.A1(_2903_),
    .A2(_2906_),
    .ZN(_2907_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _6295_ (.A1(\mod.Data_Mem.F_M.MRAM[13][4] ),
    .A2(_2901_),
    .B1(_2902_),
    .B2(\mod.Data_Mem.F_M.MRAM[12][4] ),
    .C(_2907_),
    .ZN(_2908_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6296_ (.A1(_2144_),
    .A2(\mod.Data_Mem.F_M.MRAM[783][4] ),
    .B1(\mod.Data_Mem.F_M.MRAM[782][4] ),
    .B2(_2267_),
    .ZN(_2909_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6297_ (.A1(_2752_),
    .A2(_2909_),
    .ZN(_2910_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _6298_ (.A1(\mod.Data_Mem.F_M.MRAM[781][4] ),
    .A2(_2751_),
    .B1(_2157_),
    .B2(\mod.Data_Mem.F_M.MRAM[780][4] ),
    .C(_2910_),
    .ZN(_2911_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _6299_ (.I0(_2232_),
    .I1(_2237_),
    .I2(_2908_),
    .I3(_2911_),
    .S0(_1964_),
    .S1(_2759_),
    .Z(_2912_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6300_ (.A1(_2703_),
    .A2(_2912_),
    .ZN(_2913_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6301_ (.A1(_2868_),
    .A2(_2900_),
    .B(_2913_),
    .ZN(_2914_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6302_ (.A1(_2866_),
    .A2(_2914_),
    .ZN(_0068_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6303_ (.A1(_2870_),
    .A2(_1969_),
    .ZN(_2915_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6304_ (.A1(_1664_),
    .A2(_1970_),
    .B(_2873_),
    .ZN(_2916_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6305_ (.A1(_1655_),
    .A2(_1974_),
    .ZN(_2917_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6306_ (.A1(_2876_),
    .A2(_1973_),
    .B(_2763_),
    .ZN(_2918_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6307_ (.A1(_2915_),
    .A2(_2916_),
    .B1(_2917_),
    .B2(_2918_),
    .ZN(_2919_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6308_ (.A1(_2869_),
    .A2(_2919_),
    .ZN(_2920_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6309_ (.I0(_1978_),
    .I1(_1979_),
    .S(_2723_),
    .Z(_2921_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6310_ (.I0(_1980_),
    .I1(_1981_),
    .S(_1738_),
    .Z(_2922_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _6311_ (.A1(_2882_),
    .A2(_2921_),
    .B1(_2922_),
    .B2(_2884_),
    .C(_2078_),
    .ZN(_2923_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6312_ (.A1(_2870_),
    .A2(_1950_),
    .ZN(_2924_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6313_ (.A1(_1826_),
    .A2(_1952_),
    .B(_2873_),
    .ZN(_2925_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6314_ (.A1(_2924_),
    .A2(_2925_),
    .ZN(_2926_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6315_ (.A1(_2872_),
    .A2(_1958_),
    .ZN(_2927_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6316_ (.A1(_2891_),
    .A2(_1957_),
    .ZN(_2928_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6317_ (.A1(_2718_),
    .A2(_2927_),
    .A3(_2928_),
    .ZN(_2929_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6318_ (.A1(_2886_),
    .A2(_2926_),
    .A3(_2929_),
    .ZN(_2930_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6319_ (.A1(_1603_),
    .A2(_1937_),
    .ZN(_2931_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6320_ (.A1(_1566_),
    .A2(_1936_),
    .B(_2931_),
    .ZN(_2932_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6321_ (.I0(_1943_),
    .I1(_1945_),
    .S(_2044_),
    .Z(_2933_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _6322_ (.A1(_2895_),
    .A2(_2932_),
    .B1(_2933_),
    .B2(_2898_),
    .C(_1866_),
    .ZN(_2934_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6323_ (.A1(_2920_),
    .A2(_2923_),
    .B1(_2930_),
    .B2(_2934_),
    .ZN(_2935_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6324_ (.A1(_2134_),
    .A2(\mod.Data_Mem.F_M.MRAM[15][5] ),
    .B1(\mod.Data_Mem.F_M.MRAM[14][5] ),
    .B2(_2905_),
    .ZN(_2936_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6325_ (.A1(_2903_),
    .A2(_2936_),
    .ZN(_2937_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _6326_ (.A1(\mod.Data_Mem.F_M.MRAM[13][5] ),
    .A2(_2901_),
    .B1(_2902_),
    .B2(\mod.Data_Mem.F_M.MRAM[12][5] ),
    .C(_2937_),
    .ZN(_2938_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6327_ (.A1(_2904_),
    .A2(\mod.Data_Mem.F_M.MRAM[783][5] ),
    .B1(\mod.Data_Mem.F_M.MRAM[782][5] ),
    .B2(_2267_),
    .ZN(_2939_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6328_ (.A1(_2752_),
    .A2(_2939_),
    .ZN(_2940_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _6329_ (.A1(\mod.Data_Mem.F_M.MRAM[781][5] ),
    .A2(_2751_),
    .B1(_2157_),
    .B2(\mod.Data_Mem.F_M.MRAM[780][5] ),
    .C(_2940_),
    .ZN(_2941_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _6330_ (.I0(_2240_),
    .I1(_2243_),
    .I2(_2938_),
    .I3(_2941_),
    .S0(_1964_),
    .S1(_2759_),
    .Z(_2942_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6331_ (.A1(_2867_),
    .A2(_2942_),
    .ZN(_2943_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6332_ (.A1(_2868_),
    .A2(_2935_),
    .B(_2943_),
    .ZN(_2944_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6333_ (.A1(_2866_),
    .A2(_2944_),
    .ZN(_0069_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6334_ (.A1(_2870_),
    .A2(_2004_),
    .ZN(_2945_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6335_ (.A1(_1635_),
    .A2(_2005_),
    .ZN(_2946_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6336_ (.A1(_2846_),
    .A2(_2945_),
    .A3(_2946_),
    .ZN(_2947_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6337_ (.A1(_1635_),
    .A2(_2003_),
    .ZN(_2948_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6338_ (.A1(_1941_),
    .A2(_2002_),
    .ZN(_2949_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6339_ (.A1(_2779_),
    .A2(_2948_),
    .A3(_2949_),
    .ZN(_2950_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6340_ (.A1(_2886_),
    .A2(_2947_),
    .A3(_2950_),
    .ZN(_2951_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _6341_ (.I0(\mod.Data_Mem.F_M.MRAM[789][6] ),
    .I1(\mod.Data_Mem.F_M.MRAM[791][6] ),
    .I2(\mod.Data_Mem.F_M.MRAM[790][6] ),
    .I3(\mod.Data_Mem.F_M.MRAM[788][6] ),
    .S0(_2448_),
    .S1(_1932_),
    .Z(_2952_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6342_ (.I0(_2015_),
    .I1(_2016_),
    .S(_1738_),
    .Z(_2953_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _6343_ (.A1(_2882_),
    .A2(_2952_),
    .B1(_2953_),
    .B2(_2884_),
    .C(_1898_),
    .ZN(_2954_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6344_ (.A1(_1635_),
    .A2(_1990_),
    .ZN(_2955_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6345_ (.A1(_1608_),
    .A2(_1989_),
    .B(_2763_),
    .ZN(_2956_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6346_ (.A1(_2876_),
    .A2(_1987_),
    .ZN(_2957_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6347_ (.A1(_2012_),
    .A2(_1988_),
    .B(_2739_),
    .ZN(_2958_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6348_ (.A1(_2955_),
    .A2(_2956_),
    .B1(_2957_),
    .B2(_2958_),
    .ZN(_2959_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6349_ (.A1(_2869_),
    .A2(_2959_),
    .ZN(_2960_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6350_ (.I0(_1997_),
    .I1(_1996_),
    .S(_1713_),
    .Z(_2961_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6351_ (.I0(_1994_),
    .I1(_1995_),
    .S(_2044_),
    .Z(_2962_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _6352_ (.A1(_2884_),
    .A2(_2961_),
    .B1(_2962_),
    .B2(_2895_),
    .C(_1725_),
    .ZN(_2963_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6353_ (.A1(_2951_),
    .A2(_2954_),
    .B1(_2960_),
    .B2(_2963_),
    .ZN(_2964_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6354_ (.A1(_2134_),
    .A2(\mod.Data_Mem.F_M.MRAM[15][6] ),
    .B1(\mod.Data_Mem.F_M.MRAM[14][6] ),
    .B2(_2216_),
    .ZN(_2965_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6355_ (.A1(_2903_),
    .A2(_2965_),
    .ZN(_2966_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _6356_ (.A1(\mod.Data_Mem.F_M.MRAM[13][6] ),
    .A2(_2901_),
    .B1(_2201_),
    .B2(\mod.Data_Mem.F_M.MRAM[12][6] ),
    .C(_2966_),
    .ZN(_2967_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6357_ (.A1(_2904_),
    .A2(\mod.Data_Mem.F_M.MRAM[783][6] ),
    .B1(\mod.Data_Mem.F_M.MRAM[782][6] ),
    .B2(_2905_),
    .ZN(_2968_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6358_ (.A1(_2752_),
    .A2(_2968_),
    .ZN(_2969_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _6359_ (.A1(\mod.Data_Mem.F_M.MRAM[781][6] ),
    .A2(_2751_),
    .B1(_2902_),
    .B2(\mod.Data_Mem.F_M.MRAM[780][6] ),
    .C(_2969_),
    .ZN(_2970_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _6360_ (.I0(_2246_),
    .I1(_2249_),
    .I2(_2967_),
    .I3(_2970_),
    .S0(_1964_),
    .S1(_2750_),
    .Z(_2971_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6361_ (.A1(_2867_),
    .A2(_2971_),
    .ZN(_2972_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6362_ (.A1(_2868_),
    .A2(_2964_),
    .B(_2972_),
    .ZN(_2973_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6363_ (.A1(_2866_),
    .A2(_2973_),
    .ZN(_0070_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6364_ (.A1(_1585_),
    .A2(_2026_),
    .ZN(_2974_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6365_ (.A1(_2876_),
    .A2(_2024_),
    .B(_2715_),
    .ZN(_2975_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6366_ (.A1(_1941_),
    .A2(_2027_),
    .ZN(_2976_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6367_ (.A1(_1834_),
    .A2(_2028_),
    .B(_2873_),
    .ZN(_2977_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6368_ (.A1(_2974_),
    .A2(_2975_),
    .B1(_2976_),
    .B2(_2977_),
    .ZN(_2978_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6369_ (.A1(_2869_),
    .A2(_2978_),
    .ZN(_2979_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6370_ (.I0(_2032_),
    .I1(_2033_),
    .S(_1738_),
    .Z(_2980_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6371_ (.I0(_2034_),
    .I1(_2035_),
    .S(_2180_),
    .Z(_2981_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _6372_ (.A1(_2882_),
    .A2(_2980_),
    .B1(_2981_),
    .B2(_2898_),
    .C(_2078_),
    .ZN(_2982_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6373_ (.A1(_1655_),
    .A2(_2041_),
    .ZN(_2983_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6374_ (.A1(_2891_),
    .A2(_2040_),
    .ZN(_2984_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6375_ (.A1(_2779_),
    .A2(_2983_),
    .A3(_2984_),
    .ZN(_2985_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6376_ (.A1(_2891_),
    .A2(_2042_),
    .ZN(_2986_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6377_ (.A1(_2872_),
    .A2(_2043_),
    .ZN(_2987_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6378_ (.A1(_2733_),
    .A2(_2986_),
    .A3(_2987_),
    .ZN(_2988_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6379_ (.A1(_2886_),
    .A2(_2985_),
    .A3(_2988_),
    .ZN(_2989_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _6380_ (.I0(\mod.Data_Mem.F_M.MRAM[789][7] ),
    .I1(\mod.Data_Mem.F_M.MRAM[791][7] ),
    .I2(\mod.Data_Mem.F_M.MRAM[790][7] ),
    .I3(\mod.Data_Mem.F_M.MRAM[788][7] ),
    .S0(_1915_),
    .S1(_2383_),
    .Z(_2990_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6381_ (.I0(_2051_),
    .I1(_2052_),
    .S(_1881_),
    .Z(_2991_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _6382_ (.A1(_2895_),
    .A2(_2990_),
    .B1(_2991_),
    .B2(_2898_),
    .C(_1866_),
    .ZN(_2992_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6383_ (.A1(_2979_),
    .A2(_2982_),
    .B1(_2989_),
    .B2(_2992_),
    .ZN(_2993_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6384_ (.A1(_2134_),
    .A2(\mod.Data_Mem.F_M.MRAM[15][7] ),
    .B1(\mod.Data_Mem.F_M.MRAM[14][7] ),
    .B2(_2216_),
    .ZN(_2994_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6385_ (.A1(_1565_),
    .A2(_2994_),
    .ZN(_2995_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _6386_ (.A1(\mod.Data_Mem.F_M.MRAM[13][7] ),
    .A2(_1538_),
    .B1(_2201_),
    .B2(\mod.Data_Mem.F_M.MRAM[12][7] ),
    .C(_2995_),
    .ZN(_2996_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6387_ (.A1(_2904_),
    .A2(\mod.Data_Mem.F_M.MRAM[783][7] ),
    .B1(\mod.Data_Mem.F_M.MRAM[782][7] ),
    .B2(_2905_),
    .ZN(_2997_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6388_ (.A1(_2903_),
    .A2(_2997_),
    .ZN(_2998_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _6389_ (.A1(\mod.Data_Mem.F_M.MRAM[781][7] ),
    .A2(_2901_),
    .B1(_2902_),
    .B2(\mod.Data_Mem.F_M.MRAM[780][7] ),
    .C(_2998_),
    .ZN(_2999_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _6390_ (.I0(_2252_),
    .I1(_2255_),
    .I2(_2996_),
    .I3(_2999_),
    .S0(_1489_),
    .S1(_2750_),
    .Z(_3000_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6391_ (.A1(_2867_),
    .A2(_3000_),
    .ZN(_3001_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6392_ (.A1(_2868_),
    .A2(_2993_),
    .B(_3001_),
    .ZN(_3002_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6393_ (.A1(_2866_),
    .A2(_3002_),
    .ZN(_0071_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6394_ (.I(_1724_),
    .Z(_3003_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6395_ (.I(_2698_),
    .Z(_3004_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6396_ (.I(_2092_),
    .Z(_3005_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6397_ (.I(_2429_),
    .Z(_3006_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _6398_ (.A1(_3005_),
    .A2(_2261_),
    .B1(_3006_),
    .B2(_2407_),
    .C1(_2404_),
    .C2(_2510_),
    .ZN(_3007_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6399_ (.A1(_3004_),
    .A2(_3007_),
    .ZN(_3008_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6400_ (.I(_2499_),
    .Z(_3009_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6401_ (.A1(_2418_),
    .A2(\mod.Data_Mem.F_M.MRAM[780][0] ),
    .ZN(_3010_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6402_ (.A1(_2256_),
    .A2(\mod.Data_Mem.F_M.MRAM[781][0] ),
    .ZN(_3011_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _6403_ (.A1(_2422_),
    .A2(_3010_),
    .A3(_3011_),
    .ZN(_3012_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _6404_ (.A1(_3009_),
    .A2(_2389_),
    .B1(_2384_),
    .B2(_2503_),
    .C(_3012_),
    .ZN(_3013_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6405_ (.I(_2100_),
    .Z(_3014_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _6406_ (.A1(_2110_),
    .A2(_2387_),
    .B(_3013_),
    .C(_3014_),
    .ZN(_3015_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6407_ (.A1(_3003_),
    .A2(_3008_),
    .A3(_3015_),
    .ZN(_3016_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6408_ (.I(_2385_),
    .Z(_3017_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _6409_ (.A1(_2171_),
    .A2(\mod.Data_Mem.F_M.MRAM[12][0] ),
    .Z(_3018_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _6410_ (.A1(_3017_),
    .A2(\mod.Data_Mem.F_M.MRAM[13][0] ),
    .B(_2382_),
    .C(_3018_),
    .ZN(_3019_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6411_ (.I(_2376_),
    .Z(_3020_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6412_ (.I(_3020_),
    .Z(_3021_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6413_ (.I0(\mod.Data_Mem.F_M.MRAM[0][0] ),
    .I1(\mod.Data_Mem.F_M.MRAM[1][0] ),
    .S(_2258_),
    .Z(_3022_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6414_ (.I(_2495_),
    .Z(_3023_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _6415_ (.A1(_3021_),
    .A2(_2359_),
    .B1(_3022_),
    .B2(_3023_),
    .C1(_3009_),
    .C2(_2368_),
    .ZN(_3024_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6416_ (.A1(_3014_),
    .A2(_3019_),
    .A3(_3024_),
    .ZN(_3025_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6417_ (.I(_2092_),
    .Z(_3026_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _6418_ (.A1(_3026_),
    .A2(_2272_),
    .B1(_2365_),
    .B2(_3006_),
    .C1(_2361_),
    .C2(_2672_),
    .ZN(_3027_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6419_ (.A1(_2626_),
    .A2(_3027_),
    .ZN(_3028_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6420_ (.A1(_2184_),
    .A2(_3025_),
    .A3(_3028_),
    .ZN(_3029_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6421_ (.A1(_3016_),
    .A2(_3029_),
    .ZN(_0072_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6422_ (.I(_2429_),
    .Z(_3030_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6423_ (.I(_2388_),
    .Z(_3031_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _6424_ (.A1(_2447_),
    .A2(_2278_),
    .B1(_3030_),
    .B2(_2420_),
    .C1(_2427_),
    .C2(_3031_),
    .ZN(_3032_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6425_ (.A1(_3020_),
    .A2(_2438_),
    .ZN(_3033_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _6426_ (.A1(_2301_),
    .A2(\mod.Data_Mem.F_M.MRAM[780][1] ),
    .Z(_3034_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _6427_ (.A1(_2728_),
    .A2(\mod.Data_Mem.F_M.MRAM[781][1] ),
    .B(_2381_),
    .C(_3034_),
    .ZN(_3035_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6428_ (.A1(_1933_),
    .A2(\mod.Data_Mem.F_M.MRAM[769][1] ),
    .ZN(_3036_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6429_ (.A1(_2620_),
    .A2(_1716_),
    .B(_3036_),
    .ZN(_3037_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6430_ (.A1(_2560_),
    .A2(_2437_),
    .B1(_3037_),
    .B2(_2388_),
    .ZN(_3038_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _6431_ (.A1(_1536_),
    .A2(_3033_),
    .A3(_3035_),
    .A4(_3038_),
    .ZN(_3039_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6432_ (.A1(_1965_),
    .A2(_3039_),
    .ZN(_3040_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6433_ (.A1(_2626_),
    .A2(_3032_),
    .B(_3040_),
    .ZN(_3041_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6434_ (.A1(_2343_),
    .A2(\mod.Data_Mem.F_M.MRAM[12][1] ),
    .ZN(_3042_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6435_ (.A1(_2417_),
    .A2(\mod.Data_Mem.F_M.MRAM[13][1] ),
    .ZN(_3043_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6436_ (.A1(_2071_),
    .A2(_3042_),
    .A3(_3043_),
    .ZN(_3044_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _6437_ (.A1(_2312_),
    .A2(_2459_),
    .B(_3044_),
    .C(_3026_),
    .ZN(_3045_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6438_ (.I0(\mod.Data_Mem.F_M.MRAM[0][1] ),
    .I1(\mod.Data_Mem.F_M.MRAM[1][1] ),
    .S(_2512_),
    .Z(_3046_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6439_ (.I(_1619_),
    .Z(_3047_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _6440_ (.A1(_3030_),
    .A2(_2451_),
    .B1(_3046_),
    .B2(_2672_),
    .C(_3047_),
    .ZN(_3048_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6441_ (.I(_2092_),
    .Z(_3049_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6442_ (.I(_2499_),
    .Z(_3050_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _6443_ (.A1(_3049_),
    .A2(_2285_),
    .B1(_3050_),
    .B2(_2453_),
    .C1(_2460_),
    .C2(_2496_),
    .ZN(_3051_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _6444_ (.A1(_3045_),
    .A2(_3048_),
    .B1(_3051_),
    .B2(_2831_),
    .C(_2073_),
    .ZN(_3052_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _6445_ (.A1(_3041_),
    .A2(_3052_),
    .Z(_3053_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6446_ (.I(_3053_),
    .Z(_0073_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _6447_ (.A1(_3005_),
    .A2(_2292_),
    .B1(_3006_),
    .B2(_2466_),
    .C1(_2469_),
    .C2(_3023_),
    .ZN(_3054_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6448_ (.A1(_3004_),
    .A2(_3054_),
    .ZN(_3055_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6449_ (.A1(_3017_),
    .A2(\mod.Data_Mem.F_M.MRAM[781][2] ),
    .ZN(_3056_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6450_ (.A1(_2696_),
    .A2(\mod.Data_Mem.F_M.MRAM[780][2] ),
    .B(_2382_),
    .ZN(_3057_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6451_ (.A1(_2258_),
    .A2(\mod.Data_Mem.F_M.MRAM[769][2] ),
    .ZN(_3058_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6452_ (.A1(_2345_),
    .A2(_1770_),
    .B(_3058_),
    .ZN(_3059_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6453_ (.I(_2499_),
    .Z(_3060_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _6454_ (.A1(_2503_),
    .A2(_2478_),
    .B1(_3059_),
    .B2(_2568_),
    .C1(_3060_),
    .C2(_2477_),
    .ZN(_3061_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _6455_ (.A1(_3056_),
    .A2(_3057_),
    .B(_3061_),
    .C(_3014_),
    .ZN(_3062_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6456_ (.A1(_3003_),
    .A2(_3055_),
    .A3(_3062_),
    .ZN(_3063_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6457_ (.A1(\mod.Data_Mem.F_M.MRAM[13][2] ),
    .A2(_2382_),
    .B1(_2642_),
    .B2(\mod.Data_Mem.F_M.MRAM[1][2] ),
    .ZN(_3064_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6458_ (.A1(_2063_),
    .A2(_3064_),
    .ZN(_3065_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _6459_ (.A1(_2619_),
    .A2(\mod.Data_Mem.F_M.MRAM[0][2] ),
    .Z(_3066_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _6460_ (.A1(_3021_),
    .A2(_2490_),
    .B1(_3066_),
    .B2(_3031_),
    .C(_3047_),
    .ZN(_3067_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6461_ (.A1(\mod.Data_Mem.F_M.MRAM[12][2] ),
    .A2(_1886_),
    .B1(_2536_),
    .B2(_2486_),
    .ZN(_3068_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6462_ (.A1(_3067_),
    .A2(_3068_),
    .ZN(_3069_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _6463_ (.A1(_3005_),
    .A2(_2298_),
    .B1(_3009_),
    .B2(_2487_),
    .C1(_2491_),
    .C2(_3023_),
    .ZN(_3070_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6464_ (.A1(_2831_),
    .A2(_3070_),
    .B(_2073_),
    .ZN(_3071_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6465_ (.A1(_3065_),
    .A2(_3069_),
    .B(_3071_),
    .ZN(_3072_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6466_ (.A1(_3063_),
    .A2(_3072_),
    .ZN(_0074_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _6467_ (.A1(_2171_),
    .A2(\mod.Data_Mem.F_M.MRAM[0][3] ),
    .Z(_3073_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _6468_ (.A1(_3017_),
    .A2(\mod.Data_Mem.F_M.MRAM[1][3] ),
    .B(_3031_),
    .C(_3073_),
    .ZN(_3074_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6469_ (.A1(_2151_),
    .A2(\mod.Data_Mem.F_M.MRAM[13][3] ),
    .ZN(_3075_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6470_ (.A1(_2275_),
    .A2(\mod.Data_Mem.F_M.MRAM[12][3] ),
    .ZN(_3076_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _6471_ (.A1(_2422_),
    .A2(_3075_),
    .A3(_3076_),
    .ZN(_3077_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _6472_ (.A1(_3021_),
    .A2(_2527_),
    .B1(_2524_),
    .B2(_3009_),
    .C(_3077_),
    .ZN(_3078_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6473_ (.A1(_3014_),
    .A2(_3074_),
    .A3(_3078_),
    .ZN(_3079_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _6474_ (.A1(_3026_),
    .A2(_2304_),
    .B1(_3006_),
    .B2(_2523_),
    .C1(_2529_),
    .C2(_2510_),
    .ZN(_3080_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6475_ (.A1(_3004_),
    .A2(_3080_),
    .ZN(_3081_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6476_ (.A1(_2184_),
    .A2(_3079_),
    .A3(_3081_),
    .ZN(_3082_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6477_ (.I(_2189_),
    .Z(_3083_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6478_ (.A1(_2315_),
    .A2(\mod.Data_Mem.F_M.MRAM[769][3] ),
    .ZN(_3084_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6479_ (.A1(_3083_),
    .A2(_1855_),
    .B(_3084_),
    .ZN(_3085_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6480_ (.A1(_3031_),
    .A2(_3085_),
    .B(_3047_),
    .ZN(_3086_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6481_ (.A1(_2264_),
    .A2(\mod.Data_Mem.F_M.MRAM[781][3] ),
    .ZN(_3087_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6482_ (.A1(_2475_),
    .A2(\mod.Data_Mem.F_M.MRAM[780][3] ),
    .ZN(_3088_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _6483_ (.A1(_2439_),
    .A2(_3087_),
    .A3(_3088_),
    .ZN(_3089_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6484_ (.A1(_3030_),
    .A2(_2514_),
    .B(_3089_),
    .ZN(_3090_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _6485_ (.A1(_2072_),
    .A2(_2509_),
    .B(_3086_),
    .C(_3090_),
    .ZN(_3091_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _6486_ (.A1(_3026_),
    .A2(_2309_),
    .B1(_3030_),
    .B2(_2497_),
    .C1(_2502_),
    .C2(_2672_),
    .ZN(_3092_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6487_ (.A1(_3004_),
    .A2(_3092_),
    .ZN(_3093_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6488_ (.A1(_3003_),
    .A2(_3091_),
    .A3(_3093_),
    .ZN(_3094_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6489_ (.A1(_3082_),
    .A2(_3094_),
    .ZN(_0075_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _6490_ (.I0(\mod.Data_Mem.F_M.MRAM[12][4] ),
    .I1(\mod.Data_Mem.F_M.MRAM[14][4] ),
    .I2(\mod.Data_Mem.F_M.MRAM[13][4] ),
    .I3(_1870_),
    .S0(_2290_),
    .S1(_2171_),
    .Z(_3095_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6491_ (.A1(_2728_),
    .A2(\mod.Data_Mem.F_M.MRAM[1][4] ),
    .ZN(_3096_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6492_ (.A1(_2511_),
    .A2(\mod.Data_Mem.F_M.MRAM[0][4] ),
    .B(_2103_),
    .ZN(_3097_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _6493_ (.A1(_2345_),
    .A2(\mod.Data_Mem.F_M.MRAM[2][4] ),
    .B(_2440_),
    .C(_2569_),
    .ZN(_3098_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6494_ (.A1(_3096_),
    .A2(_3097_),
    .B(_3098_),
    .ZN(_3099_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _6495_ (.A1(_2353_),
    .A2(_3095_),
    .B(_3099_),
    .C(_2108_),
    .ZN(_3100_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6496_ (.A1(_2103_),
    .A2(_2559_),
    .ZN(_3101_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6497_ (.A1(_3047_),
    .A2(_3101_),
    .ZN(_3102_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _6498_ (.A1(_2353_),
    .A2(_2318_),
    .B1(_2536_),
    .B2(_2556_),
    .C(_3102_),
    .ZN(_3103_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _6499_ (.I0(\mod.Data_Mem.F_M.MRAM[780][4] ),
    .I1(\mod.Data_Mem.F_M.MRAM[782][4] ),
    .I2(\mod.Data_Mem.F_M.MRAM[781][4] ),
    .I3(_1901_),
    .S0(_2270_),
    .S1(_3083_),
    .Z(_3104_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6500_ (.A1(_3083_),
    .A2(\mod.Data_Mem.F_M.MRAM[768][4] ),
    .ZN(_3105_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6501_ (.I(_2203_),
    .Z(_3106_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6502_ (.I(_2102_),
    .Z(_3107_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6503_ (.A1(_3106_),
    .A2(\mod.Data_Mem.F_M.MRAM[769][4] ),
    .B(_3107_),
    .ZN(_3108_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6504_ (.A1(_3105_),
    .A2(_3108_),
    .B(_2474_),
    .ZN(_3109_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _6505_ (.A1(_2611_),
    .A2(_2547_),
    .B1(_3104_),
    .B2(_2211_),
    .C(_3109_),
    .ZN(_3110_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6506_ (.I(_2107_),
    .Z(_3111_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _6507_ (.A1(_3049_),
    .A2(_2323_),
    .B1(_2500_),
    .B2(_2543_),
    .C1(_2541_),
    .C2(_2568_),
    .ZN(_3112_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6508_ (.A1(_3111_),
    .A2(_3112_),
    .ZN(_3113_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6509_ (.A1(_1491_),
    .A2(_3113_),
    .ZN(_3114_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _6510_ (.A1(_1966_),
    .A2(_3100_),
    .A3(_3103_),
    .B1(_3110_),
    .B2(_3114_),
    .ZN(_0076_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6511_ (.A1(_2587_),
    .A2(\mod.Data_Mem.F_M.MRAM[13][5] ),
    .ZN(_3115_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6512_ (.A1(_2696_),
    .A2(\mod.Data_Mem.F_M.MRAM[12][5] ),
    .B(_2596_),
    .ZN(_3116_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6513_ (.A1(_2528_),
    .A2(\mod.Data_Mem.F_M.MRAM[0][5] ),
    .ZN(_3117_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _6514_ (.A1(_2475_),
    .A2(_1971_),
    .B(_2406_),
    .C(_3117_),
    .ZN(_3118_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _6515_ (.A1(_3060_),
    .A2(_2591_),
    .B1(_2592_),
    .B2(_3020_),
    .C(_3118_),
    .ZN(_3119_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _6516_ (.A1(_3115_),
    .A2(_3116_),
    .B(_3119_),
    .C(_2434_),
    .ZN(_3120_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _6517_ (.A1(_3049_),
    .A2(_2329_),
    .B1(_3050_),
    .B2(_2578_),
    .C1(_2580_),
    .C2(_2496_),
    .ZN(_3121_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6518_ (.A1(_3111_),
    .A2(_3121_),
    .ZN(_3122_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6519_ (.A1(_3120_),
    .A2(_3122_),
    .ZN(_3123_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6520_ (.A1(_3106_),
    .A2(\mod.Data_Mem.F_M.MRAM[781][5] ),
    .ZN(_3124_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6521_ (.A1(_2567_),
    .A2(\mod.Data_Mem.F_M.MRAM[780][5] ),
    .B(_2596_),
    .ZN(_3125_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6522_ (.A1(_2321_),
    .A2(\mod.Data_Mem.F_M.MRAM[768][5] ),
    .ZN(_3126_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _6523_ (.A1(_2315_),
    .A2(_1955_),
    .B(_2406_),
    .C(_3126_),
    .ZN(_3127_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6524_ (.A1(_2500_),
    .A2(_2602_),
    .B(_3127_),
    .ZN(_3128_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _6525_ (.A1(_2558_),
    .A2(_2598_),
    .B1(_3124_),
    .B2(_3125_),
    .C(_3128_),
    .ZN(_3129_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _6526_ (.A1(_2508_),
    .A2(_2333_),
    .B1(_3060_),
    .B2(_2605_),
    .C1(_2606_),
    .C2(_3107_),
    .ZN(_3130_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6527_ (.A1(_3111_),
    .A2(_3130_),
    .ZN(_3131_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _6528_ (.A1(_2626_),
    .A2(_3129_),
    .B(_3131_),
    .C(_2079_),
    .ZN(_3132_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6529_ (.A1(_2534_),
    .A2(_3123_),
    .B(_3132_),
    .ZN(_0077_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _6530_ (.A1(_2424_),
    .A2(\mod.Data_Mem.F_M.MRAM[12][6] ),
    .Z(_3133_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _6531_ (.A1(_3106_),
    .A2(\mod.Data_Mem.F_M.MRAM[13][6] ),
    .B(_2394_),
    .C(_3133_),
    .ZN(_3134_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6532_ (.A1(_2061_),
    .A2(\mod.Data_Mem.F_M.MRAM[1][6] ),
    .ZN(_3135_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6533_ (.A1(_2522_),
    .A2(\mod.Data_Mem.F_M.MRAM[0][6] ),
    .B(_2102_),
    .ZN(_3136_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6534_ (.A1(_3135_),
    .A2(_3136_),
    .ZN(_3137_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _6535_ (.A1(_3060_),
    .A2(_2643_),
    .B1(_2644_),
    .B2(_3020_),
    .C(_3137_),
    .ZN(_3138_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _6536_ (.A1(_2474_),
    .A2(_3134_),
    .A3(_3138_),
    .Z(_3139_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _6537_ (.A1(_2071_),
    .A2(_2210_),
    .A3(_2636_),
    .B(_2698_),
    .ZN(_3140_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _6538_ (.A1(_2447_),
    .A2(_2337_),
    .B1(_2631_),
    .B2(_2642_),
    .C(_3140_),
    .ZN(_3141_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _6539_ (.A1(_2522_),
    .A2(\mod.Data_Mem.F_M.MRAM[781][6] ),
    .Z(_3142_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _6540_ (.A1(_2619_),
    .A2(\mod.Data_Mem.F_M.MRAM[780][6] ),
    .B(_3142_),
    .C(_2170_),
    .ZN(_3143_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6541_ (.A1(_2091_),
    .A2(_2622_),
    .B(_3143_),
    .ZN(_3144_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6542_ (.A1(_3083_),
    .A2(\mod.Data_Mem.F_M.MRAM[768][6] ),
    .ZN(_3145_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6543_ (.A1(_3106_),
    .A2(\mod.Data_Mem.F_M.MRAM[769][6] ),
    .B(_3107_),
    .ZN(_3146_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6544_ (.A1(_3145_),
    .A2(_3146_),
    .B(_2474_),
    .ZN(_3147_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _6545_ (.A1(_2611_),
    .A2(_2627_),
    .B1(_3144_),
    .B2(_2211_),
    .C(_3147_),
    .ZN(_3148_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _6546_ (.A1(_3049_),
    .A2(_2341_),
    .B1(_2500_),
    .B2(_2615_),
    .C1(_2616_),
    .C2(_2568_),
    .ZN(_3149_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6547_ (.A1(_3111_),
    .A2(_3149_),
    .ZN(_3150_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6548_ (.A1(_1491_),
    .A2(_3150_),
    .ZN(_3151_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _6549_ (.A1(_1966_),
    .A2(_3139_),
    .A3(_3141_),
    .B1(_3148_),
    .B2(_3151_),
    .ZN(_0078_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6550_ (.A1(_2728_),
    .A2(\mod.Data_Mem.F_M.MRAM[1][7] ),
    .ZN(_3152_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6551_ (.A1(_2511_),
    .A2(\mod.Data_Mem.F_M.MRAM[0][7] ),
    .B(_2103_),
    .ZN(_3153_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6552_ (.A1(_2417_),
    .A2(\mod.Data_Mem.F_M.MRAM[12][7] ),
    .ZN(_3154_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6553_ (.A1(_2343_),
    .A2(\mod.Data_Mem.F_M.MRAM[13][7] ),
    .B(_2381_),
    .ZN(_3155_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6554_ (.A1(_2548_),
    .A2(_2673_),
    .ZN(_3156_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _6555_ (.A1(_3152_),
    .A2(_3153_),
    .B1(_3154_),
    .B2(_3155_),
    .C(_3156_),
    .ZN(_3157_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _6556_ (.A1(_3021_),
    .A2(_2677_),
    .B(_3157_),
    .C(_2108_),
    .ZN(_3158_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _6557_ (.A1(_2312_),
    .A2(_2508_),
    .A3(_2668_),
    .B(_1757_),
    .ZN(_3159_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _6558_ (.A1(_2353_),
    .A2(_2347_),
    .B1(_2663_),
    .B2(_2642_),
    .C(_3159_),
    .ZN(_3160_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _6559_ (.A1(_3005_),
    .A2(_2350_),
    .B1(_3050_),
    .B2(_2652_),
    .C1(_2650_),
    .C2(_2496_),
    .ZN(_3161_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6560_ (.A1(_2831_),
    .A2(_3161_),
    .ZN(_3162_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6561_ (.A1(\mod.Data_Mem.F_M.MRAM[781][7] ),
    .A2(_2596_),
    .B1(_3023_),
    .B2(\mod.Data_Mem.F_M.MRAM[769][7] ),
    .ZN(_3163_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _6562_ (.A1(_2385_),
    .A2(\mod.Data_Mem.F_M.MRAM[768][7] ),
    .Z(_3164_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _6563_ (.A1(\mod.Data_Mem.F_M.MRAM[780][7] ),
    .A2(_1674_),
    .B1(_3107_),
    .B2(_3164_),
    .C(_2698_),
    .ZN(_3165_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6564_ (.A1(_2503_),
    .A2(_2655_),
    .B1(_2656_),
    .B2(_3050_),
    .ZN(_3166_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _6565_ (.A1(_3017_),
    .A2(_3163_),
    .B(_3165_),
    .C(_3166_),
    .ZN(_3167_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6566_ (.A1(_1966_),
    .A2(_3162_),
    .A3(_3167_),
    .ZN(_3168_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _6567_ (.A1(_3003_),
    .A2(_3158_),
    .A3(_3160_),
    .B(_3168_),
    .ZN(_0079_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6568_ (.I(\mod.I_addr[1] ),
    .Z(_3169_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6569_ (.A1(_0612_),
    .A2(_3169_),
    .Z(_3170_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6570_ (.I(_3170_),
    .Z(_0081_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6571_ (.I(\mod.I_addr[2] ),
    .Z(_3171_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6572_ (.A1(_0612_),
    .A2(_3169_),
    .ZN(_3172_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _6573_ (.A1(_3171_),
    .A2(_3172_),
    .ZN(_3173_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6574_ (.I(_3173_),
    .Z(_0082_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6575_ (.I(\mod.I_addr[3] ),
    .ZN(_3174_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6576_ (.I(_3174_),
    .Z(_3175_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _6577_ (.A1(\mod.I_addr[0] ),
    .A2(\mod.I_addr[2] ),
    .A3(\mod.I_addr[1] ),
    .ZN(_3176_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6578_ (.A1(_3175_),
    .A2(_3176_),
    .Z(_3177_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6579_ (.I(_3177_),
    .Z(_0083_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6580_ (.I(\mod.I_addr[4] ),
    .Z(_3178_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _6581_ (.A1(_3175_),
    .A2(_3176_),
    .ZN(_3179_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6582_ (.A1(_3178_),
    .A2(_3179_),
    .Z(_3180_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6583_ (.I(_3180_),
    .Z(_0084_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6584_ (.A1(_3178_),
    .A2(_3179_),
    .ZN(_3181_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _6585_ (.A1(\mod.I_addr[5] ),
    .A2(_3181_),
    .ZN(_3182_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6586_ (.I(_3182_),
    .Z(_0085_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6587_ (.A1(_3178_),
    .A2(\mod.I_addr[5] ),
    .A3(_3179_),
    .ZN(_3183_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _6588_ (.A1(\mod.I_addr[6] ),
    .A2(_3183_),
    .ZN(_3184_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6589_ (.I(_3184_),
    .Z(_0086_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _6590_ (.A1(_3178_),
    .A2(\mod.I_addr[6] ),
    .A3(\mod.I_addr[5] ),
    .A4(_3179_),
    .ZN(_3185_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _6591_ (.A1(\mod.I_addr[7] ),
    .A2(_3185_),
    .ZN(_3186_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6592_ (.I(_3186_),
    .Z(_0087_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6593_ (.I(\mod.Data_Mem.F_M.MRAM[11][0] ),
    .Z(_3187_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6594_ (.I(_3187_),
    .Z(_0088_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6595_ (.I(\mod.Data_Mem.F_M.MRAM[11][1] ),
    .Z(_3188_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6596_ (.I(_3188_),
    .Z(_0089_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6597_ (.I(\mod.Data_Mem.F_M.MRAM[11][2] ),
    .Z(_3189_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6598_ (.I(_3189_),
    .Z(_0090_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6599_ (.I(\mod.Data_Mem.F_M.MRAM[11][3] ),
    .Z(_3190_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6600_ (.I(_3190_),
    .Z(_0091_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6601_ (.I(\mod.Data_Mem.F_M.MRAM[11][4] ),
    .Z(_3191_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6602_ (.I(_3191_),
    .Z(_0092_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6603_ (.I(\mod.Data_Mem.F_M.MRAM[11][5] ),
    .Z(_3192_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6604_ (.I(_3192_),
    .Z(_0093_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6605_ (.I(\mod.Data_Mem.F_M.MRAM[11][6] ),
    .Z(_3193_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6606_ (.I(_3193_),
    .Z(_0094_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6607_ (.I(\mod.Data_Mem.F_M.MRAM[11][7] ),
    .Z(_3194_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6608_ (.I(_3194_),
    .Z(_0095_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6609_ (.I(\mod.Data_Mem.F_M.MRAM[24][0] ),
    .Z(_3195_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6610_ (.I(_3195_),
    .Z(_0096_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6611_ (.I(\mod.Data_Mem.F_M.MRAM[24][1] ),
    .Z(_3196_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6612_ (.I(_3196_),
    .Z(_0097_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6613_ (.I(\mod.Data_Mem.F_M.MRAM[24][2] ),
    .Z(_3197_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6614_ (.I(_3197_),
    .Z(_0098_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6615_ (.I(\mod.Data_Mem.F_M.MRAM[24][3] ),
    .Z(_3198_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6616_ (.I(_3198_),
    .Z(_0099_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6617_ (.I(\mod.Data_Mem.F_M.MRAM[24][4] ),
    .Z(_3199_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6618_ (.I(_3199_),
    .Z(_0100_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6619_ (.I(\mod.Data_Mem.F_M.MRAM[24][5] ),
    .Z(_3200_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6620_ (.I(_3200_),
    .Z(_0101_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6621_ (.I(\mod.Data_Mem.F_M.MRAM[24][6] ),
    .Z(_3201_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6622_ (.I(_3201_),
    .Z(_0102_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6623_ (.I(\mod.Data_Mem.F_M.MRAM[24][7] ),
    .Z(_3202_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6624_ (.I(_3202_),
    .Z(_0103_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6625_ (.I(\mod.Data_Mem.F_M.MRAM[26][0] ),
    .Z(_3203_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6626_ (.I(_3203_),
    .Z(_0104_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6627_ (.I(\mod.Data_Mem.F_M.MRAM[26][1] ),
    .Z(_3204_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6628_ (.I(_3204_),
    .Z(_0105_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6629_ (.I(\mod.Data_Mem.F_M.MRAM[26][2] ),
    .Z(_3205_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6630_ (.I(_3205_),
    .Z(_0106_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6631_ (.I(\mod.Data_Mem.F_M.MRAM[26][3] ),
    .Z(_3206_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6632_ (.I(_3206_),
    .Z(_0107_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6633_ (.I(\mod.Data_Mem.F_M.MRAM[26][4] ),
    .Z(_3207_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6634_ (.I(_3207_),
    .Z(_0108_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6635_ (.I(\mod.Data_Mem.F_M.MRAM[26][5] ),
    .Z(_3208_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6636_ (.I(_3208_),
    .Z(_0109_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6637_ (.I(\mod.Data_Mem.F_M.MRAM[26][6] ),
    .Z(_3209_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6638_ (.I(_3209_),
    .Z(_0110_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6639_ (.I(\mod.Data_Mem.F_M.MRAM[26][7] ),
    .Z(_3210_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6640_ (.I(_3210_),
    .Z(_0111_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6641_ (.I(\mod.Data_Mem.F_M.MRAM[25][0] ),
    .Z(_3211_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6642_ (.I(_3211_),
    .Z(_0112_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6643_ (.I(\mod.Data_Mem.F_M.MRAM[25][1] ),
    .Z(_3212_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6644_ (.I(_3212_),
    .Z(_0113_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6645_ (.I(\mod.Data_Mem.F_M.MRAM[25][2] ),
    .Z(_3213_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6646_ (.I(_3213_),
    .Z(_0114_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6647_ (.I(\mod.Data_Mem.F_M.MRAM[25][3] ),
    .Z(_3214_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6648_ (.I(_3214_),
    .Z(_0115_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6649_ (.I(\mod.Data_Mem.F_M.MRAM[25][4] ),
    .Z(_3215_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6650_ (.I(_3215_),
    .Z(_0116_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6651_ (.I(\mod.Data_Mem.F_M.MRAM[25][5] ),
    .Z(_3216_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6652_ (.I(_3216_),
    .Z(_0117_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6653_ (.I(\mod.Data_Mem.F_M.MRAM[25][6] ),
    .Z(_3217_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6654_ (.I(_3217_),
    .Z(_0118_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6655_ (.I(\mod.Data_Mem.F_M.MRAM[25][7] ),
    .Z(_3218_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6656_ (.I(_3218_),
    .Z(_0119_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6657_ (.I(\mod.Data_Mem.F_M.MRAM[27][0] ),
    .Z(_3219_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6658_ (.I(_3219_),
    .Z(_0120_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6659_ (.I(\mod.Data_Mem.F_M.MRAM[27][1] ),
    .Z(_3220_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6660_ (.I(_3220_),
    .Z(_0121_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6661_ (.I(\mod.Data_Mem.F_M.MRAM[27][2] ),
    .Z(_3221_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6662_ (.I(_3221_),
    .Z(_0122_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6663_ (.I(\mod.Data_Mem.F_M.MRAM[27][3] ),
    .Z(_3222_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6664_ (.I(_3222_),
    .Z(_0123_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6665_ (.I(\mod.Data_Mem.F_M.MRAM[27][4] ),
    .Z(_3223_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6666_ (.I(_3223_),
    .Z(_0124_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6667_ (.I(\mod.Data_Mem.F_M.MRAM[27][5] ),
    .Z(_3224_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6668_ (.I(_3224_),
    .Z(_0125_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6669_ (.I(\mod.Data_Mem.F_M.MRAM[27][6] ),
    .Z(_3225_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6670_ (.I(_3225_),
    .Z(_0126_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6671_ (.I(\mod.Data_Mem.F_M.MRAM[27][7] ),
    .Z(_3226_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6672_ (.I(_3226_),
    .Z(_0127_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6673_ (.I(net3),
    .Z(_3227_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6674_ (.I(_3227_),
    .Z(_3228_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _6675_ (.A1(\mod.Data_Mem.F_M.dest[4] ),
    .A2(\mod.Data_Mem.F_M.dest[2] ),
    .Z(_3229_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6676_ (.I(_3229_),
    .Z(_3230_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6677_ (.A1(\mod.Data_Mem.F_M.dest[1] ),
    .A2(\mod.Data_Mem.F_M.dest[0] ),
    .ZN(_3231_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6678_ (.I(_3231_),
    .Z(_3232_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6679_ (.I(\mod.DMen_reg2 ),
    .ZN(_3233_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6680_ (.A1(\mod.Data_Mem.F_M.dest[8] ),
    .A2(_3233_),
    .ZN(_3234_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6681_ (.I(_3234_),
    .Z(_3235_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6682_ (.A1(_3230_),
    .A2(_3232_),
    .A3(_3235_),
    .ZN(_3236_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _6683_ (.I(_3236_),
    .Z(_3237_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6684_ (.I0(_3228_),
    .I1(\mod.Data_Mem.F_M.MRAM[28][0] ),
    .S(_3237_),
    .Z(_3238_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6685_ (.I(_3238_),
    .Z(_0128_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6686_ (.I(net4),
    .Z(_3239_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6687_ (.I(_3239_),
    .Z(_3240_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6688_ (.I0(_3240_),
    .I1(\mod.Data_Mem.F_M.MRAM[28][1] ),
    .S(_3237_),
    .Z(_3241_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6689_ (.I(_3241_),
    .Z(_0129_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6690_ (.I(net5),
    .Z(_3242_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6691_ (.I(_3242_),
    .Z(_3243_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6692_ (.I0(_3243_),
    .I1(\mod.Data_Mem.F_M.MRAM[28][2] ),
    .S(_3237_),
    .Z(_3244_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6693_ (.I(_3244_),
    .Z(_0130_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6694_ (.I(net6),
    .Z(_3245_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6695_ (.I(_3245_),
    .Z(_3246_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6696_ (.I0(_3246_),
    .I1(\mod.Data_Mem.F_M.MRAM[28][3] ),
    .S(_3237_),
    .Z(_3247_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6697_ (.I(_3247_),
    .Z(_0131_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6698_ (.I(net7),
    .Z(_3248_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6699_ (.I(_3248_),
    .Z(_3249_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _6700_ (.I(_3236_),
    .Z(_3250_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6701_ (.I0(_3249_),
    .I1(\mod.Data_Mem.F_M.MRAM[28][4] ),
    .S(_3250_),
    .Z(_3251_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6702_ (.I(_3251_),
    .Z(_0132_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6703_ (.I(net8),
    .Z(_3252_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6704_ (.I(_3252_),
    .Z(_3253_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6705_ (.I0(_3253_),
    .I1(\mod.Data_Mem.F_M.MRAM[28][5] ),
    .S(_3250_),
    .Z(_3254_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6706_ (.I(_3254_),
    .Z(_0133_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6707_ (.I(net9),
    .Z(_3255_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6708_ (.I(_3255_),
    .Z(_3256_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6709_ (.I0(_3256_),
    .I1(\mod.Data_Mem.F_M.MRAM[28][6] ),
    .S(_3250_),
    .Z(_3257_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6710_ (.I(_3257_),
    .Z(_0134_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6711_ (.I(net10),
    .Z(_3258_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6712_ (.I(_3258_),
    .Z(_3259_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6713_ (.I0(_3259_),
    .I1(\mod.Data_Mem.F_M.MRAM[28][7] ),
    .S(_3250_),
    .Z(_3260_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6714_ (.I(_3260_),
    .Z(_0135_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6715_ (.I(\mod.Data_Mem.F_M.MRAM[10][0] ),
    .Z(_3261_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6716_ (.I(_3261_),
    .Z(_0136_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6717_ (.I(\mod.Data_Mem.F_M.MRAM[10][1] ),
    .Z(_3262_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6718_ (.I(_3262_),
    .Z(_0137_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6719_ (.I(\mod.Data_Mem.F_M.MRAM[10][2] ),
    .Z(_3263_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6720_ (.I(_3263_),
    .Z(_0138_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6721_ (.I(\mod.Data_Mem.F_M.MRAM[10][3] ),
    .Z(_3264_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6722_ (.I(_3264_),
    .Z(_0139_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6723_ (.I(\mod.Data_Mem.F_M.MRAM[10][4] ),
    .Z(_3265_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6724_ (.I(_3265_),
    .Z(_0140_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6725_ (.I(\mod.Data_Mem.F_M.MRAM[10][5] ),
    .Z(_3266_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6726_ (.I(_3266_),
    .Z(_0141_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6727_ (.I(\mod.Data_Mem.F_M.MRAM[10][6] ),
    .Z(_3267_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6728_ (.I(_3267_),
    .Z(_0142_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6729_ (.I(\mod.Data_Mem.F_M.MRAM[10][7] ),
    .Z(_3268_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6730_ (.I(_3268_),
    .Z(_0143_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6731_ (.I(_3231_),
    .Z(_3269_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6732_ (.I(_3234_),
    .Z(_3270_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6733_ (.A1(\mod.Data_Mem.F_M.dest[4] ),
    .A2(\mod.Data_Mem.F_M.dest[2] ),
    .ZN(_3271_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6734_ (.I(_3271_),
    .Z(_3272_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6735_ (.A1(_3269_),
    .A2(_3270_),
    .A3(_3272_),
    .ZN(_3273_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _6736_ (.I(_3273_),
    .Z(_3274_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6737_ (.I0(_3228_),
    .I1(\mod.Data_Mem.F_M.MRAM[0][0] ),
    .S(_3274_),
    .Z(_3275_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6738_ (.I(_3275_),
    .Z(_0144_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6739_ (.I0(_3240_),
    .I1(\mod.Data_Mem.F_M.MRAM[0][1] ),
    .S(_3274_),
    .Z(_3276_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6740_ (.I(_3276_),
    .Z(_0145_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6741_ (.I0(_3243_),
    .I1(\mod.Data_Mem.F_M.MRAM[0][2] ),
    .S(_3274_),
    .Z(_3277_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6742_ (.I(_3277_),
    .Z(_0146_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6743_ (.I0(_3246_),
    .I1(\mod.Data_Mem.F_M.MRAM[0][3] ),
    .S(_3274_),
    .Z(_3278_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6744_ (.I(_3278_),
    .Z(_0147_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _6745_ (.I(_3273_),
    .Z(_3279_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6746_ (.I0(_3249_),
    .I1(\mod.Data_Mem.F_M.MRAM[0][4] ),
    .S(_3279_),
    .Z(_3280_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6747_ (.I(_3280_),
    .Z(_0148_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6748_ (.I0(_3253_),
    .I1(\mod.Data_Mem.F_M.MRAM[0][5] ),
    .S(_3279_),
    .Z(_3281_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6749_ (.I(_3281_),
    .Z(_0149_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6750_ (.I0(_3256_),
    .I1(\mod.Data_Mem.F_M.MRAM[0][6] ),
    .S(_3279_),
    .Z(_3282_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6751_ (.I(_3282_),
    .Z(_0150_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6752_ (.I0(_3259_),
    .I1(\mod.Data_Mem.F_M.MRAM[0][7] ),
    .S(_3279_),
    .Z(_3283_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6753_ (.I(_3283_),
    .Z(_0151_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6754_ (.I(\mod.Data_Mem.F_M.MRAM[8][0] ),
    .Z(_3284_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6755_ (.I(_3284_),
    .Z(_0152_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6756_ (.I(\mod.Data_Mem.F_M.MRAM[8][1] ),
    .Z(_3285_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6757_ (.I(_3285_),
    .Z(_0153_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6758_ (.I(\mod.Data_Mem.F_M.MRAM[8][2] ),
    .Z(_3286_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6759_ (.I(_3286_),
    .Z(_0154_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6760_ (.I(\mod.Data_Mem.F_M.MRAM[8][3] ),
    .Z(_3287_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6761_ (.I(_3287_),
    .Z(_0155_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6762_ (.I(\mod.Data_Mem.F_M.MRAM[8][4] ),
    .Z(_3288_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6763_ (.I(_3288_),
    .Z(_0156_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6764_ (.I(\mod.Data_Mem.F_M.MRAM[8][5] ),
    .Z(_3289_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6765_ (.I(_3289_),
    .Z(_0157_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6766_ (.I(\mod.Data_Mem.F_M.MRAM[8][6] ),
    .Z(_3290_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6767_ (.I(_3290_),
    .Z(_0158_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6768_ (.I(\mod.Data_Mem.F_M.MRAM[8][7] ),
    .Z(_3291_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6769_ (.I(_3291_),
    .Z(_0159_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6770_ (.I(net3),
    .Z(_3292_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6771_ (.I(_3292_),
    .Z(_3293_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6772_ (.I(_3229_),
    .Z(_3294_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _6773_ (.A1(\mod.Data_Mem.F_M.dest[1] ),
    .A2(\mod.Data_Mem.F_M.dest[0] ),
    .Z(_3295_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6774_ (.I(_3295_),
    .Z(_3296_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _6775_ (.A1(\mod.Data_Mem.F_M.dest[8] ),
    .A2(\mod.DMen_reg2 ),
    .Z(_3297_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6776_ (.I(_3297_),
    .Z(_3298_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _6777_ (.A1(_3294_),
    .A2(_3296_),
    .A3(_3298_),
    .Z(_3299_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _6778_ (.I(_3299_),
    .Z(_3300_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6779_ (.I0(\mod.Data_Mem.F_M.MRAM[799][0] ),
    .I1(_3293_),
    .S(_3300_),
    .Z(_3301_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6780_ (.I(_3301_),
    .Z(_0160_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6781_ (.I(net4),
    .Z(_3302_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6782_ (.I(_3302_),
    .Z(_3303_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6783_ (.I0(\mod.Data_Mem.F_M.MRAM[799][1] ),
    .I1(_3303_),
    .S(_3300_),
    .Z(_3304_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6784_ (.I(_3304_),
    .Z(_0161_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6785_ (.I(net5),
    .Z(_3305_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6786_ (.I(_3305_),
    .Z(_3306_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6787_ (.I0(\mod.Data_Mem.F_M.MRAM[799][2] ),
    .I1(_3306_),
    .S(_3300_),
    .Z(_3307_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6788_ (.I(_3307_),
    .Z(_0162_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6789_ (.I(net6),
    .Z(_3308_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6790_ (.I(_3308_),
    .Z(_3309_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6791_ (.I0(\mod.Data_Mem.F_M.MRAM[799][3] ),
    .I1(_3309_),
    .S(_3300_),
    .Z(_3310_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6792_ (.I(_3310_),
    .Z(_0163_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6793_ (.I(net7),
    .Z(_3311_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6794_ (.I(_3311_),
    .Z(_3312_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _6795_ (.I(_3299_),
    .Z(_3313_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6796_ (.I0(\mod.Data_Mem.F_M.MRAM[799][4] ),
    .I1(_3312_),
    .S(_3313_),
    .Z(_3314_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6797_ (.I(_3314_),
    .Z(_0164_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6798_ (.I(net8),
    .Z(_3315_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6799_ (.I(_3315_),
    .Z(_3316_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6800_ (.I0(\mod.Data_Mem.F_M.MRAM[799][5] ),
    .I1(_3316_),
    .S(_3313_),
    .Z(_3317_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6801_ (.I(_3317_),
    .Z(_0165_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6802_ (.I(net9),
    .Z(_3318_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6803_ (.I(_3318_),
    .Z(_3319_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6804_ (.I0(\mod.Data_Mem.F_M.MRAM[799][6] ),
    .I1(_3319_),
    .S(_3313_),
    .Z(_3320_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6805_ (.I(_3320_),
    .Z(_0166_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6806_ (.I(net10),
    .Z(_3321_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6807_ (.I(_3321_),
    .Z(_3322_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6808_ (.I0(\mod.Data_Mem.F_M.MRAM[799][7] ),
    .I1(_3322_),
    .S(_3313_),
    .Z(_3323_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6809_ (.I(_3323_),
    .Z(_0167_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6810_ (.I(\mod.Data_Mem.F_M.MRAM[789][0] ),
    .Z(_3324_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6811_ (.I(_3324_),
    .Z(_0168_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6812_ (.I(\mod.Data_Mem.F_M.MRAM[789][1] ),
    .Z(_3325_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6813_ (.I(_3325_),
    .Z(_0169_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6814_ (.I(\mod.Data_Mem.F_M.MRAM[789][2] ),
    .Z(_3326_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6815_ (.I(_3326_),
    .Z(_0170_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6816_ (.I(\mod.Data_Mem.F_M.MRAM[789][3] ),
    .Z(_3327_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6817_ (.I(_3327_),
    .Z(_0171_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6818_ (.I(\mod.Data_Mem.F_M.MRAM[789][4] ),
    .Z(_3328_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6819_ (.I(_3328_),
    .Z(_0172_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6820_ (.I(\mod.Data_Mem.F_M.MRAM[789][5] ),
    .Z(_3329_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6821_ (.I(_3329_),
    .Z(_0173_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6822_ (.I(\mod.Data_Mem.F_M.MRAM[789][6] ),
    .Z(_3330_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6823_ (.I(_3330_),
    .Z(_0174_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6824_ (.I(\mod.Data_Mem.F_M.MRAM[789][7] ),
    .Z(_3331_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6825_ (.I(_3331_),
    .Z(_0175_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6826_ (.I(_3271_),
    .Z(_3332_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6827_ (.I(\mod.Data_Mem.F_M.dest[0] ),
    .ZN(_3333_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6828_ (.A1(\mod.Data_Mem.F_M.dest[1] ),
    .A2(_3333_),
    .ZN(_3334_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _6829_ (.I(_3334_),
    .Z(_3335_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _6830_ (.A1(_3332_),
    .A2(_3298_),
    .A3(_3335_),
    .ZN(_3336_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _6831_ (.I(_3336_),
    .Z(_3337_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6832_ (.I0(_3228_),
    .I1(\mod.Data_Mem.F_M.MRAM[769][0] ),
    .S(_3337_),
    .Z(_3338_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6833_ (.I(_3338_),
    .Z(_0176_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6834_ (.I0(_3240_),
    .I1(\mod.Data_Mem.F_M.MRAM[769][1] ),
    .S(_3337_),
    .Z(_3339_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6835_ (.I(_3339_),
    .Z(_0177_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _6836_ (.I(_3336_),
    .Z(_3340_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6837_ (.I0(_3243_),
    .I1(\mod.Data_Mem.F_M.MRAM[769][2] ),
    .S(_3340_),
    .Z(_3341_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6838_ (.I(_3341_),
    .Z(_0178_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6839_ (.I0(_3246_),
    .I1(\mod.Data_Mem.F_M.MRAM[769][3] ),
    .S(_3340_),
    .Z(_3342_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6840_ (.I(_3342_),
    .Z(_0179_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6841_ (.I0(_3249_),
    .I1(\mod.Data_Mem.F_M.MRAM[769][4] ),
    .S(_3340_),
    .Z(_3343_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6842_ (.I(_3343_),
    .Z(_0180_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6843_ (.A1(_3316_),
    .A2(_3337_),
    .ZN(_3344_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6844_ (.A1(_1955_),
    .A2(_3337_),
    .B(_3344_),
    .ZN(_0181_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6845_ (.I0(_3256_),
    .I1(\mod.Data_Mem.F_M.MRAM[769][6] ),
    .S(_3340_),
    .Z(_3345_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6846_ (.I(_3345_),
    .Z(_0182_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6847_ (.I0(_3259_),
    .I1(\mod.Data_Mem.F_M.MRAM[769][7] ),
    .S(_3336_),
    .Z(_3346_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6848_ (.I(_3346_),
    .Z(_0183_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6849_ (.I(\mod.Data_Mem.F_M.MRAM[779][0] ),
    .Z(_3347_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6850_ (.I(_3347_),
    .Z(_0184_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6851_ (.I(\mod.Data_Mem.F_M.MRAM[779][1] ),
    .Z(_3348_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6852_ (.I(_3348_),
    .Z(_0185_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6853_ (.I(\mod.Data_Mem.F_M.MRAM[779][2] ),
    .Z(_3349_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6854_ (.I(_3349_),
    .Z(_0186_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6855_ (.I(\mod.Data_Mem.F_M.MRAM[779][3] ),
    .Z(_3350_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6856_ (.I(_3350_),
    .Z(_0187_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6857_ (.I(\mod.Data_Mem.F_M.MRAM[779][4] ),
    .Z(_3351_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6858_ (.I(_3351_),
    .Z(_0188_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6859_ (.I(\mod.Data_Mem.F_M.MRAM[779][5] ),
    .Z(_3352_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6860_ (.I(_3352_),
    .Z(_0189_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6861_ (.I(\mod.Data_Mem.F_M.MRAM[779][6] ),
    .Z(_3353_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6862_ (.I(_3353_),
    .Z(_0190_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6863_ (.I(\mod.Data_Mem.F_M.MRAM[779][7] ),
    .Z(_3354_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6864_ (.I(_3354_),
    .Z(_0191_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6865_ (.I(\mod.Data_Mem.F_M.MRAM[6][0] ),
    .Z(_3355_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6866_ (.I(_3355_),
    .Z(_0192_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6867_ (.I(\mod.Data_Mem.F_M.MRAM[6][1] ),
    .Z(_3356_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6868_ (.I(_3356_),
    .Z(_0193_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6869_ (.I(\mod.Data_Mem.F_M.MRAM[6][2] ),
    .Z(_3357_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6870_ (.I(_3357_),
    .Z(_0194_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6871_ (.I(\mod.Data_Mem.F_M.MRAM[6][3] ),
    .Z(_3358_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6872_ (.I(_3358_),
    .Z(_0195_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6873_ (.I(\mod.Data_Mem.F_M.MRAM[6][4] ),
    .Z(_3359_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6874_ (.I(_3359_),
    .Z(_0196_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6875_ (.I(\mod.Data_Mem.F_M.MRAM[6][5] ),
    .Z(_3360_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6876_ (.I(_3360_),
    .Z(_0197_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6877_ (.I(\mod.Data_Mem.F_M.MRAM[6][6] ),
    .Z(_3361_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6878_ (.I(_3361_),
    .Z(_0198_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6879_ (.I(\mod.Data_Mem.F_M.MRAM[6][7] ),
    .Z(_3362_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6880_ (.I(_3362_),
    .Z(_0199_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6881_ (.I(\mod.Data_Mem.F_M.MRAM[4][0] ),
    .Z(_3363_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6882_ (.I(_3363_),
    .Z(_0200_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6883_ (.I(\mod.Data_Mem.F_M.MRAM[4][1] ),
    .Z(_3364_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6884_ (.I(_3364_),
    .Z(_0201_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6885_ (.I(\mod.Data_Mem.F_M.MRAM[4][2] ),
    .Z(_3365_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6886_ (.I(_3365_),
    .Z(_0202_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6887_ (.I(\mod.Data_Mem.F_M.MRAM[4][3] ),
    .Z(_3366_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6888_ (.I(_3366_),
    .Z(_0203_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6889_ (.I(\mod.Data_Mem.F_M.MRAM[4][4] ),
    .Z(_3367_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6890_ (.I(_3367_),
    .Z(_0204_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6891_ (.I(\mod.Data_Mem.F_M.MRAM[4][5] ),
    .Z(_3368_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6892_ (.I(_3368_),
    .Z(_0205_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6893_ (.I(\mod.Data_Mem.F_M.MRAM[4][6] ),
    .Z(_3369_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6894_ (.I(_3369_),
    .Z(_0206_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6895_ (.I(\mod.Data_Mem.F_M.MRAM[4][7] ),
    .Z(_3370_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6896_ (.I(_3370_),
    .Z(_0207_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6897_ (.I(_3334_),
    .Z(_3371_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6898_ (.I(\mod.Data_Mem.F_M.dest[2] ),
    .ZN(_3372_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6899_ (.A1(\mod.Data_Mem.F_M.dest[4] ),
    .A2(_3372_),
    .ZN(_3373_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6900_ (.I(_3373_),
    .Z(_3374_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6901_ (.A1(_3235_),
    .A2(_3371_),
    .A3(_3374_),
    .ZN(_3375_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _6902_ (.I(_3375_),
    .Z(_3376_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6903_ (.I0(_3228_),
    .I1(\mod.Data_Mem.F_M.MRAM[13][0] ),
    .S(_3376_),
    .Z(_3377_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6904_ (.I(_3377_),
    .Z(_0208_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6905_ (.I0(_3240_),
    .I1(\mod.Data_Mem.F_M.MRAM[13][1] ),
    .S(_3376_),
    .Z(_3378_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6906_ (.I(_3378_),
    .Z(_0209_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6907_ (.I0(_3243_),
    .I1(\mod.Data_Mem.F_M.MRAM[13][2] ),
    .S(_3376_),
    .Z(_3379_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6908_ (.I(_3379_),
    .Z(_0210_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6909_ (.I0(_3246_),
    .I1(\mod.Data_Mem.F_M.MRAM[13][3] ),
    .S(_3376_),
    .Z(_3380_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6910_ (.I(_3380_),
    .Z(_0211_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _6911_ (.I(_3375_),
    .Z(_3381_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6912_ (.I0(_3249_),
    .I1(\mod.Data_Mem.F_M.MRAM[13][4] ),
    .S(_3381_),
    .Z(_3382_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6913_ (.I(_3382_),
    .Z(_0212_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6914_ (.I0(_3253_),
    .I1(\mod.Data_Mem.F_M.MRAM[13][5] ),
    .S(_3381_),
    .Z(_3383_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6915_ (.I(_3383_),
    .Z(_0213_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6916_ (.I0(_3256_),
    .I1(\mod.Data_Mem.F_M.MRAM[13][6] ),
    .S(_3381_),
    .Z(_3384_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6917_ (.I(_3384_),
    .Z(_0214_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6918_ (.I0(_3259_),
    .I1(\mod.Data_Mem.F_M.MRAM[13][7] ),
    .S(_3381_),
    .Z(_3385_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6919_ (.I(_3385_),
    .Z(_0215_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6920_ (.I(_3227_),
    .Z(_3386_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6921_ (.I(_3373_),
    .Z(_3387_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _6922_ (.A1(\mod.Data_Mem.F_M.dest[1] ),
    .A2(_3333_),
    .Z(_3388_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6923_ (.I(_3388_),
    .Z(_3389_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6924_ (.A1(_3235_),
    .A2(_3387_),
    .A3(_3389_),
    .ZN(_3390_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _6925_ (.I(_3390_),
    .Z(_3391_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6926_ (.I0(_3386_),
    .I1(\mod.Data_Mem.F_M.MRAM[14][0] ),
    .S(_3391_),
    .Z(_3392_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6927_ (.I(_3392_),
    .Z(_0216_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6928_ (.I(_3239_),
    .Z(_3393_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6929_ (.I0(_3393_),
    .I1(\mod.Data_Mem.F_M.MRAM[14][1] ),
    .S(_3391_),
    .Z(_3394_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6930_ (.I(_3394_),
    .Z(_0217_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6931_ (.I(_3242_),
    .Z(_3395_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6932_ (.I0(_3395_),
    .I1(\mod.Data_Mem.F_M.MRAM[14][2] ),
    .S(_3391_),
    .Z(_3396_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6933_ (.I(_3396_),
    .Z(_0218_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6934_ (.I(_3245_),
    .Z(_3397_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6935_ (.I0(_3397_),
    .I1(\mod.Data_Mem.F_M.MRAM[14][3] ),
    .S(_3391_),
    .Z(_3398_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6936_ (.I(_3398_),
    .Z(_0219_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6937_ (.I(_3248_),
    .Z(_3399_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _6938_ (.I(_3390_),
    .Z(_3400_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6939_ (.I0(_3399_),
    .I1(\mod.Data_Mem.F_M.MRAM[14][4] ),
    .S(_3400_),
    .Z(_3401_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6940_ (.I(_3401_),
    .Z(_0220_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6941_ (.I0(_3253_),
    .I1(\mod.Data_Mem.F_M.MRAM[14][5] ),
    .S(_3400_),
    .Z(_3402_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6942_ (.I(_3402_),
    .Z(_0221_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6943_ (.I(_3255_),
    .Z(_3403_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6944_ (.I0(_3403_),
    .I1(\mod.Data_Mem.F_M.MRAM[14][6] ),
    .S(_3400_),
    .Z(_3404_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6945_ (.I(_3404_),
    .Z(_0222_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6946_ (.I(_3258_),
    .Z(_3405_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6947_ (.I0(_3405_),
    .I1(\mod.Data_Mem.F_M.MRAM[14][7] ),
    .S(_3400_),
    .Z(_3406_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6948_ (.I(_3406_),
    .Z(_0223_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6949_ (.I(_3295_),
    .Z(_3407_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6950_ (.A1(_3235_),
    .A2(_3407_),
    .A3(_3374_),
    .ZN(_3408_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _6951_ (.I(_3408_),
    .Z(_3409_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6952_ (.I0(_3386_),
    .I1(\mod.Data_Mem.F_M.MRAM[15][0] ),
    .S(_3409_),
    .Z(_3410_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6953_ (.I(_3410_),
    .Z(_0224_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6954_ (.I0(_3393_),
    .I1(\mod.Data_Mem.F_M.MRAM[15][1] ),
    .S(_3409_),
    .Z(_3411_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6955_ (.I(_3411_),
    .Z(_0225_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6956_ (.I0(_3395_),
    .I1(\mod.Data_Mem.F_M.MRAM[15][2] ),
    .S(_3409_),
    .Z(_3412_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6957_ (.I(_3412_),
    .Z(_0226_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6958_ (.I0(_3397_),
    .I1(\mod.Data_Mem.F_M.MRAM[15][3] ),
    .S(_3409_),
    .Z(_3413_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6959_ (.I(_3413_),
    .Z(_0227_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _6960_ (.I(_3408_),
    .Z(_3414_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6961_ (.I0(_3399_),
    .I1(_1870_),
    .S(_3414_),
    .Z(_3415_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6962_ (.I(_3415_),
    .Z(_0228_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6963_ (.I(_3252_),
    .Z(_3416_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6964_ (.I0(_3416_),
    .I1(\mod.Data_Mem.F_M.MRAM[15][5] ),
    .S(_3414_),
    .Z(_3417_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6965_ (.I(_3417_),
    .Z(_0229_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6966_ (.I0(_3403_),
    .I1(\mod.Data_Mem.F_M.MRAM[15][6] ),
    .S(_3414_),
    .Z(_3418_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6967_ (.I(_3418_),
    .Z(_0230_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6968_ (.I0(_3405_),
    .I1(\mod.Data_Mem.F_M.MRAM[15][7] ),
    .S(_3414_),
    .Z(_3419_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6969_ (.I(_3419_),
    .Z(_0231_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _6970_ (.A1(\mod.Data_Mem.F_M.dest[4] ),
    .A2(_3372_),
    .Z(_3420_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6971_ (.I(_3420_),
    .Z(_3421_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6972_ (.A1(_3269_),
    .A2(_3270_),
    .A3(_3421_),
    .ZN(_3422_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _6973_ (.I(_3422_),
    .Z(_3423_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6974_ (.I0(_3386_),
    .I1(\mod.Data_Mem.F_M.MRAM[16][0] ),
    .S(_3423_),
    .Z(_3424_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6975_ (.I(_3424_),
    .Z(_0232_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6976_ (.I0(_3393_),
    .I1(\mod.Data_Mem.F_M.MRAM[16][1] ),
    .S(_3423_),
    .Z(_3425_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6977_ (.I(_3425_),
    .Z(_0233_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6978_ (.I0(_3395_),
    .I1(\mod.Data_Mem.F_M.MRAM[16][2] ),
    .S(_3423_),
    .Z(_3426_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6979_ (.I(_3426_),
    .Z(_0234_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6980_ (.I0(_3397_),
    .I1(\mod.Data_Mem.F_M.MRAM[16][3] ),
    .S(_3423_),
    .Z(_3427_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6981_ (.I(_3427_),
    .Z(_0235_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _6982_ (.I(_3422_),
    .Z(_3428_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6983_ (.I0(_3399_),
    .I1(\mod.Data_Mem.F_M.MRAM[16][4] ),
    .S(_3428_),
    .Z(_3429_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6984_ (.I(_3429_),
    .Z(_0236_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6985_ (.I0(_3416_),
    .I1(\mod.Data_Mem.F_M.MRAM[16][5] ),
    .S(_3428_),
    .Z(_3430_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6986_ (.I(_3430_),
    .Z(_0237_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6987_ (.I0(_3403_),
    .I1(\mod.Data_Mem.F_M.MRAM[16][6] ),
    .S(_3428_),
    .Z(_3431_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6988_ (.I(_3431_),
    .Z(_0238_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6989_ (.I0(_3405_),
    .I1(\mod.Data_Mem.F_M.MRAM[16][7] ),
    .S(_3428_),
    .Z(_3432_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6990_ (.I(_3432_),
    .Z(_0239_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6991_ (.I(_3234_),
    .Z(_3433_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6992_ (.A1(_3433_),
    .A2(_3371_),
    .A3(_3421_),
    .ZN(_3434_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _6993_ (.I(_3434_),
    .Z(_3435_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6994_ (.I0(_3386_),
    .I1(\mod.Data_Mem.F_M.MRAM[17][0] ),
    .S(_3435_),
    .Z(_3436_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6995_ (.I(_3436_),
    .Z(_0240_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6996_ (.I0(_3393_),
    .I1(\mod.Data_Mem.F_M.MRAM[17][1] ),
    .S(_3435_),
    .Z(_3437_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6997_ (.I(_3437_),
    .Z(_0241_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6998_ (.I0(_3395_),
    .I1(\mod.Data_Mem.F_M.MRAM[17][2] ),
    .S(_3435_),
    .Z(_3438_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6999_ (.I(_3438_),
    .Z(_0242_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _7000_ (.I0(_3397_),
    .I1(\mod.Data_Mem.F_M.MRAM[17][3] ),
    .S(_3435_),
    .Z(_3439_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7001_ (.I(_3439_),
    .Z(_0243_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _7002_ (.I(_3434_),
    .Z(_3440_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _7003_ (.I0(_3399_),
    .I1(\mod.Data_Mem.F_M.MRAM[17][4] ),
    .S(_3440_),
    .Z(_3441_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7004_ (.I(_3441_),
    .Z(_0244_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _7005_ (.I0(_3416_),
    .I1(\mod.Data_Mem.F_M.MRAM[17][5] ),
    .S(_3440_),
    .Z(_3442_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7006_ (.I(_3442_),
    .Z(_0245_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _7007_ (.I0(_3403_),
    .I1(\mod.Data_Mem.F_M.MRAM[17][6] ),
    .S(_3440_),
    .Z(_3443_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7008_ (.I(_3443_),
    .Z(_0246_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _7009_ (.I0(_3405_),
    .I1(\mod.Data_Mem.F_M.MRAM[17][7] ),
    .S(_3440_),
    .Z(_3444_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7010_ (.I(_3444_),
    .Z(_0247_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7011_ (.I(_3227_),
    .Z(_3445_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _7012_ (.I(_3388_),
    .Z(_3446_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _7013_ (.A1(_3433_),
    .A2(_3446_),
    .A3(_3421_),
    .ZN(_3447_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _7014_ (.I(_3447_),
    .Z(_3448_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _7015_ (.I0(_3445_),
    .I1(\mod.Data_Mem.F_M.MRAM[18][0] ),
    .S(_3448_),
    .Z(_3449_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7016_ (.I(_3449_),
    .Z(_0248_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7017_ (.I(_3239_),
    .Z(_3450_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _7018_ (.I0(_3450_),
    .I1(\mod.Data_Mem.F_M.MRAM[18][1] ),
    .S(_3448_),
    .Z(_3451_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7019_ (.I(_3451_),
    .Z(_0249_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7020_ (.I(_3242_),
    .Z(_3452_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _7021_ (.I0(_3452_),
    .I1(\mod.Data_Mem.F_M.MRAM[18][2] ),
    .S(_3448_),
    .Z(_3453_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7022_ (.I(_3453_),
    .Z(_0250_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7023_ (.I(_3245_),
    .Z(_3454_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _7024_ (.I0(_3454_),
    .I1(\mod.Data_Mem.F_M.MRAM[18][3] ),
    .S(_3448_),
    .Z(_3455_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7025_ (.I(_3455_),
    .Z(_0251_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7026_ (.I(_3248_),
    .Z(_3456_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _7027_ (.I(_3447_),
    .Z(_3457_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _7028_ (.I0(_3456_),
    .I1(\mod.Data_Mem.F_M.MRAM[18][4] ),
    .S(_3457_),
    .Z(_3458_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7029_ (.I(_3458_),
    .Z(_0252_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _7030_ (.I0(_3416_),
    .I1(\mod.Data_Mem.F_M.MRAM[18][5] ),
    .S(_3457_),
    .Z(_3459_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7031_ (.I(_3459_),
    .Z(_0253_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7032_ (.I(_3255_),
    .Z(_3460_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _7033_ (.I0(_3460_),
    .I1(\mod.Data_Mem.F_M.MRAM[18][6] ),
    .S(_3457_),
    .Z(_3461_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7034_ (.I(_3461_),
    .Z(_0254_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7035_ (.I(_3258_),
    .Z(_3462_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _7036_ (.I0(_3462_),
    .I1(\mod.Data_Mem.F_M.MRAM[18][7] ),
    .S(_3457_),
    .Z(_3463_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7037_ (.I(_3463_),
    .Z(_0255_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7038_ (.I(_3234_),
    .Z(_3464_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _7039_ (.A1(_3464_),
    .A2(_3332_),
    .A3(_3335_),
    .ZN(_3465_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _7040_ (.I(_3465_),
    .Z(_3466_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _7041_ (.I0(_3445_),
    .I1(\mod.Data_Mem.F_M.MRAM[1][0] ),
    .S(_3466_),
    .Z(_3467_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7042_ (.I(_3467_),
    .Z(_0256_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _7043_ (.I0(_3450_),
    .I1(\mod.Data_Mem.F_M.MRAM[1][1] ),
    .S(_3466_),
    .Z(_3468_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7044_ (.I(_3468_),
    .Z(_0257_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _7045_ (.I(_3465_),
    .Z(_3469_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _7046_ (.I0(_3452_),
    .I1(\mod.Data_Mem.F_M.MRAM[1][2] ),
    .S(_3469_),
    .Z(_3470_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7047_ (.I(_3470_),
    .Z(_0258_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _7048_ (.I0(_3454_),
    .I1(\mod.Data_Mem.F_M.MRAM[1][3] ),
    .S(_3469_),
    .Z(_3471_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7049_ (.I(_3471_),
    .Z(_0259_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _7050_ (.I0(_3456_),
    .I1(\mod.Data_Mem.F_M.MRAM[1][4] ),
    .S(_3469_),
    .Z(_3472_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7051_ (.I(_3472_),
    .Z(_0260_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7052_ (.A1(_3316_),
    .A2(_3466_),
    .ZN(_3473_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7053_ (.A1(_1971_),
    .A2(_3466_),
    .B(_3473_),
    .ZN(_0261_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _7054_ (.I0(_3460_),
    .I1(\mod.Data_Mem.F_M.MRAM[1][6] ),
    .S(_3469_),
    .Z(_3474_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7055_ (.I(_3474_),
    .Z(_0262_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _7056_ (.I0(_3462_),
    .I1(\mod.Data_Mem.F_M.MRAM[1][7] ),
    .S(_3465_),
    .Z(_3475_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7057_ (.I(_3475_),
    .Z(_0263_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7058_ (.I(\mod.Data_Mem.F_M.MRAM[20][0] ),
    .Z(_3476_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7059_ (.I(_3476_),
    .Z(_0264_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7060_ (.I(\mod.Data_Mem.F_M.MRAM[20][1] ),
    .Z(_3477_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7061_ (.I(_3477_),
    .Z(_0265_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7062_ (.I(\mod.Data_Mem.F_M.MRAM[20][2] ),
    .Z(_3478_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7063_ (.I(_3478_),
    .Z(_0266_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7064_ (.I(\mod.Data_Mem.F_M.MRAM[20][3] ),
    .Z(_3479_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7065_ (.I(_3479_),
    .Z(_0267_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7066_ (.I(\mod.Data_Mem.F_M.MRAM[20][4] ),
    .Z(_3480_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7067_ (.I(_3480_),
    .Z(_0268_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7068_ (.I(\mod.Data_Mem.F_M.MRAM[20][5] ),
    .Z(_3481_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7069_ (.I(_3481_),
    .Z(_0269_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7070_ (.I(\mod.Data_Mem.F_M.MRAM[20][6] ),
    .Z(_3482_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7071_ (.I(_3482_),
    .Z(_0270_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7072_ (.I(\mod.Data_Mem.F_M.MRAM[20][7] ),
    .Z(_3483_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7073_ (.I(_3483_),
    .Z(_0271_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7074_ (.I(\mod.Data_Mem.F_M.MRAM[21][0] ),
    .Z(_3484_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7075_ (.I(_3484_),
    .Z(_0272_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7076_ (.I(\mod.Data_Mem.F_M.MRAM[21][1] ),
    .Z(_3485_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7077_ (.I(_3485_),
    .Z(_0273_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7078_ (.I(\mod.Data_Mem.F_M.MRAM[21][2] ),
    .Z(_3486_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7079_ (.I(_3486_),
    .Z(_0274_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7080_ (.I(\mod.Data_Mem.F_M.MRAM[21][3] ),
    .Z(_3487_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7081_ (.I(_3487_),
    .Z(_0275_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7082_ (.I(\mod.Data_Mem.F_M.MRAM[21][4] ),
    .Z(_3488_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7083_ (.I(_3488_),
    .Z(_0276_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7084_ (.I(\mod.Data_Mem.F_M.MRAM[21][5] ),
    .Z(_3489_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7085_ (.I(_3489_),
    .Z(_0277_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7086_ (.I(\mod.Data_Mem.F_M.MRAM[21][6] ),
    .Z(_3490_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7087_ (.I(_3490_),
    .Z(_0278_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7088_ (.I(\mod.Data_Mem.F_M.MRAM[21][7] ),
    .Z(_3491_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7089_ (.I(_3491_),
    .Z(_0279_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7090_ (.I(\mod.Data_Mem.F_M.MRAM[23][0] ),
    .Z(_3492_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7091_ (.I(_3492_),
    .Z(_0280_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7092_ (.I(\mod.Data_Mem.F_M.MRAM[23][1] ),
    .Z(_3493_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7093_ (.I(_3493_),
    .Z(_0281_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7094_ (.I(\mod.Data_Mem.F_M.MRAM[23][2] ),
    .Z(_3494_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7095_ (.I(_3494_),
    .Z(_0282_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7096_ (.I(\mod.Data_Mem.F_M.MRAM[23][3] ),
    .Z(_3495_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7097_ (.I(_3495_),
    .Z(_0283_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7098_ (.I(\mod.Data_Mem.F_M.MRAM[23][4] ),
    .Z(_3496_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7099_ (.I(_3496_),
    .Z(_0284_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7100_ (.I(\mod.Data_Mem.F_M.MRAM[23][5] ),
    .Z(_3497_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7101_ (.I(_3497_),
    .Z(_0285_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7102_ (.I(\mod.Data_Mem.F_M.MRAM[23][6] ),
    .Z(_3498_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7103_ (.I(_3498_),
    .Z(_0286_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7104_ (.I(\mod.Data_Mem.F_M.MRAM[23][7] ),
    .Z(_3499_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7105_ (.I(_3499_),
    .Z(_0287_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _7106_ (.A1(_3433_),
    .A2(_3272_),
    .A3(_3407_),
    .ZN(_3500_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _7107_ (.I(_3500_),
    .Z(_3501_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _7108_ (.I0(_3445_),
    .I1(\mod.Data_Mem.F_M.MRAM[3][0] ),
    .S(_3501_),
    .Z(_3502_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7109_ (.I(_3502_),
    .Z(_0288_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _7110_ (.I0(_3450_),
    .I1(\mod.Data_Mem.F_M.MRAM[3][1] ),
    .S(_3501_),
    .Z(_3503_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7111_ (.I(_3503_),
    .Z(_0289_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _7112_ (.I0(_3452_),
    .I1(\mod.Data_Mem.F_M.MRAM[3][2] ),
    .S(_3501_),
    .Z(_3504_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7113_ (.I(_3504_),
    .Z(_0290_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _7114_ (.I0(_3454_),
    .I1(\mod.Data_Mem.F_M.MRAM[3][3] ),
    .S(_3501_),
    .Z(_3505_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7115_ (.I(_3505_),
    .Z(_0291_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _7116_ (.I(_3500_),
    .Z(_3506_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _7117_ (.I0(_3456_),
    .I1(\mod.Data_Mem.F_M.MRAM[3][4] ),
    .S(_3506_),
    .Z(_3507_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7118_ (.I(_3507_),
    .Z(_0292_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7119_ (.I(_3252_),
    .Z(_3508_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _7120_ (.I0(_3508_),
    .I1(\mod.Data_Mem.F_M.MRAM[3][5] ),
    .S(_3506_),
    .Z(_3509_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7121_ (.I(_3509_),
    .Z(_0293_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _7122_ (.I0(_3460_),
    .I1(\mod.Data_Mem.F_M.MRAM[3][6] ),
    .S(_3506_),
    .Z(_3510_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7123_ (.I(_3510_),
    .Z(_0294_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _7124_ (.I0(_3462_),
    .I1(\mod.Data_Mem.F_M.MRAM[3][7] ),
    .S(_3506_),
    .Z(_3511_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7125_ (.I(_3511_),
    .Z(_0295_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _7126_ (.A1(_3433_),
    .A2(_3407_),
    .A3(_3421_),
    .ZN(_3512_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _7127_ (.I(_3512_),
    .Z(_3513_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _7128_ (.I0(_3445_),
    .I1(\mod.Data_Mem.F_M.MRAM[19][0] ),
    .S(_3513_),
    .Z(_3514_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7129_ (.I(_3514_),
    .Z(_0296_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _7130_ (.I0(_3450_),
    .I1(\mod.Data_Mem.F_M.MRAM[19][1] ),
    .S(_3513_),
    .Z(_3515_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7131_ (.I(_3515_),
    .Z(_0297_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _7132_ (.I0(_3452_),
    .I1(\mod.Data_Mem.F_M.MRAM[19][2] ),
    .S(_3513_),
    .Z(_3516_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7133_ (.I(_3516_),
    .Z(_0298_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _7134_ (.I0(_3454_),
    .I1(\mod.Data_Mem.F_M.MRAM[19][3] ),
    .S(_3513_),
    .Z(_3517_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7135_ (.I(_3517_),
    .Z(_0299_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _7136_ (.I(_3512_),
    .Z(_3518_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _7137_ (.I0(_3456_),
    .I1(\mod.Data_Mem.F_M.MRAM[19][4] ),
    .S(_3518_),
    .Z(_3519_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7138_ (.I(_3519_),
    .Z(_0300_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _7139_ (.I0(_3508_),
    .I1(\mod.Data_Mem.F_M.MRAM[19][5] ),
    .S(_3518_),
    .Z(_3520_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7140_ (.I(_3520_),
    .Z(_0301_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _7141_ (.I0(_3460_),
    .I1(\mod.Data_Mem.F_M.MRAM[19][6] ),
    .S(_3518_),
    .Z(_3521_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7142_ (.I(_3521_),
    .Z(_0302_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _7143_ (.I0(_3462_),
    .I1(\mod.Data_Mem.F_M.MRAM[19][7] ),
    .S(_3518_),
    .Z(_3522_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7144_ (.I(_3522_),
    .Z(_0303_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7145_ (.I(_3227_),
    .Z(_3523_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _7146_ (.A1(_3269_),
    .A2(_3270_),
    .A3(_3374_),
    .ZN(_3524_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _7147_ (.I(_3524_),
    .Z(_3525_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _7148_ (.I0(_3523_),
    .I1(\mod.Data_Mem.F_M.MRAM[12][0] ),
    .S(_3525_),
    .Z(_3526_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7149_ (.I(_3526_),
    .Z(_0304_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7150_ (.I(_3239_),
    .Z(_3527_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _7151_ (.I0(_3527_),
    .I1(\mod.Data_Mem.F_M.MRAM[12][1] ),
    .S(_3525_),
    .Z(_3528_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7152_ (.I(_3528_),
    .Z(_0305_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7153_ (.I(_3242_),
    .Z(_3529_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _7154_ (.I0(_3529_),
    .I1(\mod.Data_Mem.F_M.MRAM[12][2] ),
    .S(_3525_),
    .Z(_3530_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7155_ (.I(_3530_),
    .Z(_0306_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7156_ (.I(_3245_),
    .Z(_3531_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _7157_ (.I0(_3531_),
    .I1(\mod.Data_Mem.F_M.MRAM[12][3] ),
    .S(_3525_),
    .Z(_3532_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7158_ (.I(_3532_),
    .Z(_0307_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7159_ (.I(_3248_),
    .Z(_3533_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _7160_ (.I(_3524_),
    .Z(_3534_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _7161_ (.I0(_3533_),
    .I1(\mod.Data_Mem.F_M.MRAM[12][4] ),
    .S(_3534_),
    .Z(_3535_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7162_ (.I(_3535_),
    .Z(_0308_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _7163_ (.I0(_3508_),
    .I1(\mod.Data_Mem.F_M.MRAM[12][5] ),
    .S(_3534_),
    .Z(_3536_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7164_ (.I(_3536_),
    .Z(_0309_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7165_ (.I(_3255_),
    .Z(_3537_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _7166_ (.I0(_3537_),
    .I1(\mod.Data_Mem.F_M.MRAM[12][6] ),
    .S(_3534_),
    .Z(_3538_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7167_ (.I(_3538_),
    .Z(_0310_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7168_ (.I(_3258_),
    .Z(_3539_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _7169_ (.I0(_3539_),
    .I1(\mod.Data_Mem.F_M.MRAM[12][7] ),
    .S(_3534_),
    .Z(_3540_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7170_ (.I(_3540_),
    .Z(_0311_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7171_ (.I(\mod.Data_Mem.F_M.MRAM[22][0] ),
    .Z(_3541_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7172_ (.I(_3541_),
    .Z(_0312_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7173_ (.I(\mod.Data_Mem.F_M.MRAM[22][1] ),
    .Z(_3542_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7174_ (.I(_3542_),
    .Z(_0313_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7175_ (.I(\mod.Data_Mem.F_M.MRAM[22][2] ),
    .Z(_3543_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7176_ (.I(_3543_),
    .Z(_0314_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7177_ (.I(\mod.Data_Mem.F_M.MRAM[22][3] ),
    .Z(_3544_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7178_ (.I(_3544_),
    .Z(_0315_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7179_ (.I(\mod.Data_Mem.F_M.MRAM[22][4] ),
    .Z(_3545_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7180_ (.I(_3545_),
    .Z(_0316_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7181_ (.I(\mod.Data_Mem.F_M.MRAM[22][5] ),
    .Z(_3546_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7182_ (.I(_3546_),
    .Z(_0317_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7183_ (.I(\mod.Data_Mem.F_M.MRAM[22][6] ),
    .Z(_3547_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7184_ (.I(_3547_),
    .Z(_0318_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7185_ (.I(\mod.Data_Mem.F_M.MRAM[22][7] ),
    .Z(_3548_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7186_ (.I(_3548_),
    .Z(_0319_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _7187_ (.A1(_3294_),
    .A2(_3464_),
    .A3(_3335_),
    .ZN(_3549_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _7188_ (.I(_3549_),
    .Z(_3550_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _7189_ (.I0(_3523_),
    .I1(\mod.Data_Mem.F_M.MRAM[29][0] ),
    .S(_3550_),
    .Z(_3551_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7190_ (.I(_3551_),
    .Z(_0320_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _7191_ (.I0(_3527_),
    .I1(\mod.Data_Mem.F_M.MRAM[29][1] ),
    .S(_3550_),
    .Z(_3552_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7192_ (.I(_3552_),
    .Z(_0321_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _7193_ (.I(_3549_),
    .Z(_3553_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _7194_ (.I0(_3529_),
    .I1(\mod.Data_Mem.F_M.MRAM[29][2] ),
    .S(_3553_),
    .Z(_3554_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7195_ (.I(_3554_),
    .Z(_0322_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7196_ (.I(_3308_),
    .Z(_3555_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7197_ (.A1(_3555_),
    .A2(_3550_),
    .ZN(_3556_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7198_ (.A1(_2213_),
    .A2(_3550_),
    .B(_3556_),
    .ZN(_0323_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _7199_ (.I0(_3533_),
    .I1(\mod.Data_Mem.F_M.MRAM[29][4] ),
    .S(_3553_),
    .Z(_3557_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7200_ (.I(_3557_),
    .Z(_0324_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _7201_ (.I0(_3508_),
    .I1(\mod.Data_Mem.F_M.MRAM[29][5] ),
    .S(_3553_),
    .Z(_3558_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7202_ (.I(_3558_),
    .Z(_0325_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _7203_ (.I0(_3537_),
    .I1(\mod.Data_Mem.F_M.MRAM[29][6] ),
    .S(_3553_),
    .Z(_3559_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7204_ (.I(_3559_),
    .Z(_0326_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _7205_ (.I0(_3539_),
    .I1(\mod.Data_Mem.F_M.MRAM[29][7] ),
    .S(_3549_),
    .Z(_3560_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7206_ (.I(_3560_),
    .Z(_0327_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _7207_ (.A1(_3270_),
    .A2(_3272_),
    .A3(_3389_),
    .ZN(_3561_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _7208_ (.I(_3561_),
    .Z(_3562_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _7209_ (.I0(_3523_),
    .I1(\mod.Data_Mem.F_M.MRAM[2][0] ),
    .S(_3562_),
    .Z(_3563_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7210_ (.I(_3563_),
    .Z(_0328_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _7211_ (.I0(_3527_),
    .I1(\mod.Data_Mem.F_M.MRAM[2][1] ),
    .S(_3562_),
    .Z(_3564_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7212_ (.I(_3564_),
    .Z(_0329_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _7213_ (.I0(_3529_),
    .I1(\mod.Data_Mem.F_M.MRAM[2][2] ),
    .S(_3562_),
    .Z(_3565_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7214_ (.I(_3565_),
    .Z(_0330_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _7215_ (.I0(_3531_),
    .I1(\mod.Data_Mem.F_M.MRAM[2][3] ),
    .S(_3562_),
    .Z(_3566_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7216_ (.I(_3566_),
    .Z(_0331_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _7217_ (.I(_3561_),
    .Z(_3567_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _7218_ (.I0(_3533_),
    .I1(\mod.Data_Mem.F_M.MRAM[2][4] ),
    .S(_3567_),
    .Z(_3568_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7219_ (.I(_3568_),
    .Z(_0332_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7220_ (.I(_3252_),
    .Z(_3569_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _7221_ (.I0(_3569_),
    .I1(\mod.Data_Mem.F_M.MRAM[2][5] ),
    .S(_3567_),
    .Z(_3570_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7222_ (.I(_3570_),
    .Z(_0333_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _7223_ (.I0(_3537_),
    .I1(\mod.Data_Mem.F_M.MRAM[2][6] ),
    .S(_3567_),
    .Z(_3571_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7224_ (.I(_3571_),
    .Z(_0334_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _7225_ (.I0(_3539_),
    .I1(\mod.Data_Mem.F_M.MRAM[2][7] ),
    .S(_3567_),
    .Z(_3572_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7226_ (.I(_3572_),
    .Z(_0335_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _7227_ (.A1(_3230_),
    .A2(_3464_),
    .A3(_3389_),
    .ZN(_3573_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _7228_ (.I(_3573_),
    .Z(_3574_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _7229_ (.I0(_3523_),
    .I1(\mod.Data_Mem.F_M.MRAM[30][0] ),
    .S(_3574_),
    .Z(_3575_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7230_ (.I(_3575_),
    .Z(_0336_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _7231_ (.I0(_3527_),
    .I1(\mod.Data_Mem.F_M.MRAM[30][1] ),
    .S(_3574_),
    .Z(_3576_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7232_ (.I(_3576_),
    .Z(_0337_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _7233_ (.I0(_3529_),
    .I1(\mod.Data_Mem.F_M.MRAM[30][2] ),
    .S(_3574_),
    .Z(_3577_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7234_ (.I(_3577_),
    .Z(_0338_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _7235_ (.I0(_3531_),
    .I1(\mod.Data_Mem.F_M.MRAM[30][3] ),
    .S(_3574_),
    .Z(_3578_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7236_ (.I(_3578_),
    .Z(_0339_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _7237_ (.I(_3573_),
    .Z(_3579_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _7238_ (.I0(_3533_),
    .I1(\mod.Data_Mem.F_M.MRAM[30][4] ),
    .S(_3579_),
    .Z(_3580_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7239_ (.I(_3580_),
    .Z(_0340_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _7240_ (.I0(_3569_),
    .I1(\mod.Data_Mem.F_M.MRAM[30][5] ),
    .S(_3579_),
    .Z(_3581_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7241_ (.I(_3581_),
    .Z(_0341_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _7242_ (.I0(_3537_),
    .I1(\mod.Data_Mem.F_M.MRAM[30][6] ),
    .S(_3579_),
    .Z(_3582_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7243_ (.I(_3582_),
    .Z(_0342_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _7244_ (.I0(_3539_),
    .I1(\mod.Data_Mem.F_M.MRAM[30][7] ),
    .S(_3579_),
    .Z(_3583_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7245_ (.I(_3583_),
    .Z(_0343_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _7246_ (.A1(_3294_),
    .A2(_3464_),
    .A3(_3296_),
    .Z(_3584_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _7247_ (.I(_3584_),
    .Z(_3585_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _7248_ (.I0(\mod.Data_Mem.F_M.MRAM[31][0] ),
    .I1(_3293_),
    .S(_3585_),
    .Z(_3586_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7249_ (.I(_3586_),
    .Z(_0344_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _7250_ (.I0(_1632_),
    .I1(_3303_),
    .S(_3585_),
    .Z(_3587_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7251_ (.I(_3587_),
    .Z(_0345_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _7252_ (.I0(\mod.Data_Mem.F_M.MRAM[31][2] ),
    .I1(_3306_),
    .S(_3585_),
    .Z(_3588_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7253_ (.I(_3588_),
    .Z(_0346_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _7254_ (.I0(\mod.Data_Mem.F_M.MRAM[31][3] ),
    .I1(_3555_),
    .S(_3585_),
    .Z(_3589_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7255_ (.I(_3589_),
    .Z(_0347_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _7256_ (.I(_3584_),
    .Z(_3590_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _7257_ (.I0(\mod.Data_Mem.F_M.MRAM[31][4] ),
    .I1(_3312_),
    .S(_3590_),
    .Z(_3591_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7258_ (.I(_3591_),
    .Z(_0348_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _7259_ (.I0(\mod.Data_Mem.F_M.MRAM[31][5] ),
    .I1(_3316_),
    .S(_3590_),
    .Z(_3592_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7260_ (.I(_3592_),
    .Z(_0349_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _7261_ (.I0(\mod.Data_Mem.F_M.MRAM[31][6] ),
    .I1(_3319_),
    .S(_3590_),
    .Z(_3593_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7262_ (.I(_3593_),
    .Z(_0350_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _7263_ (.I0(\mod.Data_Mem.F_M.MRAM[31][7] ),
    .I1(_3322_),
    .S(_3590_),
    .Z(_3594_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7264_ (.I(_3594_),
    .Z(_0351_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7265_ (.I(\mod.Data_Mem.F_M.MRAM[5][0] ),
    .Z(_3595_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7266_ (.I(_3595_),
    .Z(_0352_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7267_ (.I(\mod.Data_Mem.F_M.MRAM[5][1] ),
    .Z(_3596_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7268_ (.I(_3596_),
    .Z(_0353_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7269_ (.I(\mod.Data_Mem.F_M.MRAM[5][2] ),
    .Z(_3597_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7270_ (.I(_3597_),
    .Z(_0354_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7271_ (.I(\mod.Data_Mem.F_M.MRAM[5][3] ),
    .Z(_3598_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7272_ (.I(_3598_),
    .Z(_0355_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7273_ (.I(\mod.Data_Mem.F_M.MRAM[5][4] ),
    .Z(_3599_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7274_ (.I(_3599_),
    .Z(_0356_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7275_ (.I(\mod.Data_Mem.F_M.MRAM[5][5] ),
    .Z(_3600_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7276_ (.I(_3600_),
    .Z(_0357_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7277_ (.I(\mod.Data_Mem.F_M.MRAM[5][6] ),
    .Z(_3601_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7278_ (.I(_3601_),
    .Z(_0358_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7279_ (.I(\mod.Data_Mem.F_M.MRAM[5][7] ),
    .Z(_3602_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7280_ (.I(_3602_),
    .Z(_0359_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7281_ (.I(_3292_),
    .Z(_3603_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7282_ (.I(_3297_),
    .Z(_3604_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _7283_ (.A1(_3232_),
    .A2(_3332_),
    .A3(_3604_),
    .ZN(_3605_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _7284_ (.I(_3605_),
    .Z(_3606_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _7285_ (.I0(_3603_),
    .I1(\mod.Data_Mem.F_M.MRAM[768][0] ),
    .S(_3606_),
    .Z(_3607_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7286_ (.I(_3607_),
    .Z(_0360_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _7287_ (.I(_3605_),
    .Z(_3608_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7288_ (.I(_3608_),
    .Z(_3609_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7289_ (.I(_3302_),
    .Z(_3610_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7290_ (.A1(_3610_),
    .A2(_3609_),
    .ZN(_3611_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7291_ (.A1(_1716_),
    .A2(_3609_),
    .B(_3611_),
    .ZN(_0361_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7292_ (.I(_3305_),
    .Z(_3612_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7293_ (.A1(_3612_),
    .A2(_3606_),
    .ZN(_3613_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7294_ (.A1(_1770_),
    .A2(_3609_),
    .B(_3613_),
    .ZN(_0362_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7295_ (.A1(_3555_),
    .A2(_3606_),
    .ZN(_3614_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7296_ (.A1(_1855_),
    .A2(_3609_),
    .B(_3614_),
    .ZN(_0363_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7297_ (.I(_3311_),
    .Z(_3615_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _7298_ (.I0(_3615_),
    .I1(\mod.Data_Mem.F_M.MRAM[768][4] ),
    .S(_3606_),
    .Z(_3616_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7299_ (.I(_3616_),
    .Z(_0364_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _7300_ (.I0(_3569_),
    .I1(\mod.Data_Mem.F_M.MRAM[768][5] ),
    .S(_3608_),
    .Z(_3617_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7301_ (.I(_3617_),
    .Z(_0365_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7302_ (.I(_3318_),
    .Z(_3618_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _7303_ (.I0(_3618_),
    .I1(\mod.Data_Mem.F_M.MRAM[768][6] ),
    .S(_3608_),
    .Z(_3619_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7304_ (.I(_3619_),
    .Z(_0366_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7305_ (.I(_3321_),
    .Z(_3620_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _7306_ (.I0(_3620_),
    .I1(\mod.Data_Mem.F_M.MRAM[768][7] ),
    .S(_3608_),
    .Z(_3621_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7307_ (.I(_3621_),
    .Z(_0367_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _7308_ (.A1(_3332_),
    .A2(_3604_),
    .A3(_3446_),
    .ZN(_3622_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _7309_ (.I(_3622_),
    .Z(_3623_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _7310_ (.I0(_3603_),
    .I1(\mod.Data_Mem.F_M.MRAM[770][0] ),
    .S(_3623_),
    .Z(_3624_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7311_ (.I(_3624_),
    .Z(_0368_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _7312_ (.I(_3622_),
    .Z(_3625_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7313_ (.I(_3625_),
    .Z(_3626_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7314_ (.A1(_3610_),
    .A2(_3626_),
    .ZN(_3627_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7315_ (.A1(_1709_),
    .A2(_3626_),
    .B(_3627_),
    .ZN(_0369_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7316_ (.A1(_3612_),
    .A2(_3623_),
    .ZN(_3628_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7317_ (.A1(_1765_),
    .A2(_3626_),
    .B(_3628_),
    .ZN(_0370_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7318_ (.A1(_3555_),
    .A2(_3623_),
    .ZN(_3629_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7319_ (.A1(_1851_),
    .A2(_3626_),
    .B(_3629_),
    .ZN(_0371_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _7320_ (.I0(_3615_),
    .I1(\mod.Data_Mem.F_M.MRAM[770][4] ),
    .S(_3623_),
    .Z(_3630_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7321_ (.I(_3630_),
    .Z(_0372_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _7322_ (.I0(_3569_),
    .I1(\mod.Data_Mem.F_M.MRAM[770][5] ),
    .S(_3625_),
    .Z(_3631_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7323_ (.I(_3631_),
    .Z(_0373_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _7324_ (.I0(_3618_),
    .I1(\mod.Data_Mem.F_M.MRAM[770][6] ),
    .S(_3625_),
    .Z(_3632_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7325_ (.I(_3632_),
    .Z(_0374_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _7326_ (.I0(_3620_),
    .I1(\mod.Data_Mem.F_M.MRAM[770][7] ),
    .S(_3625_),
    .Z(_3633_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7327_ (.I(_3633_),
    .Z(_0375_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7328_ (.I(_3297_),
    .Z(_3634_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _7329_ (.A1(_3272_),
    .A2(_3296_),
    .A3(_3634_),
    .ZN(_3635_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _7330_ (.I(_3635_),
    .Z(_3636_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _7331_ (.I0(_3603_),
    .I1(\mod.Data_Mem.F_M.MRAM[771][0] ),
    .S(_3636_),
    .Z(_3637_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7332_ (.I(_3637_),
    .Z(_0376_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7333_ (.I(_3302_),
    .Z(_3638_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _7334_ (.I0(_3638_),
    .I1(\mod.Data_Mem.F_M.MRAM[771][1] ),
    .S(_3636_),
    .Z(_3639_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7335_ (.I(_3639_),
    .Z(_0377_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7336_ (.I(_3305_),
    .Z(_3640_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _7337_ (.I0(_3640_),
    .I1(\mod.Data_Mem.F_M.MRAM[771][2] ),
    .S(_3636_),
    .Z(_3641_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7338_ (.I(_3641_),
    .Z(_0378_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _7339_ (.I0(_3531_),
    .I1(\mod.Data_Mem.F_M.MRAM[771][3] ),
    .S(_3636_),
    .Z(_3642_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7340_ (.I(_3642_),
    .Z(_0379_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _7341_ (.I(_3635_),
    .Z(_3643_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _7342_ (.I0(_3615_),
    .I1(\mod.Data_Mem.F_M.MRAM[771][4] ),
    .S(_3643_),
    .Z(_3644_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7343_ (.I(_3644_),
    .Z(_0380_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7344_ (.I(_3315_),
    .Z(_3645_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _7345_ (.I0(_3645_),
    .I1(\mod.Data_Mem.F_M.MRAM[771][5] ),
    .S(_3643_),
    .Z(_3646_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7346_ (.I(_3646_),
    .Z(_0381_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _7347_ (.I0(_3618_),
    .I1(\mod.Data_Mem.F_M.MRAM[771][6] ),
    .S(_3643_),
    .Z(_3647_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7348_ (.I(_3647_),
    .Z(_0382_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _7349_ (.I0(_3620_),
    .I1(\mod.Data_Mem.F_M.MRAM[771][7] ),
    .S(_3643_),
    .Z(_3648_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7350_ (.I(_3648_),
    .Z(_0383_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7351_ (.I(\mod.Data_Mem.F_M.MRAM[772][0] ),
    .Z(_3649_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7352_ (.I(_3649_),
    .Z(_0384_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7353_ (.I(\mod.Data_Mem.F_M.MRAM[772][1] ),
    .Z(_3650_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7354_ (.I(_3650_),
    .Z(_0385_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7355_ (.I(\mod.Data_Mem.F_M.MRAM[772][2] ),
    .Z(_3651_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7356_ (.I(_3651_),
    .Z(_0386_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7357_ (.I(\mod.Data_Mem.F_M.MRAM[772][3] ),
    .Z(_3652_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7358_ (.I(_3652_),
    .Z(_0387_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7359_ (.I(\mod.Data_Mem.F_M.MRAM[772][4] ),
    .Z(_3653_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7360_ (.I(_3653_),
    .Z(_0388_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7361_ (.I(\mod.Data_Mem.F_M.MRAM[772][5] ),
    .Z(_3654_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7362_ (.I(_3654_),
    .Z(_0389_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7363_ (.I(\mod.Data_Mem.F_M.MRAM[772][6] ),
    .Z(_3655_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7364_ (.I(_3655_),
    .Z(_0390_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7365_ (.I(\mod.Data_Mem.F_M.MRAM[772][7] ),
    .Z(_3656_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7366_ (.I(_3656_),
    .Z(_0391_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7367_ (.I(\mod.Data_Mem.F_M.MRAM[773][0] ),
    .Z(_3657_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7368_ (.I(_3657_),
    .Z(_0392_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7369_ (.I(\mod.Data_Mem.F_M.MRAM[773][1] ),
    .Z(_3658_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7370_ (.I(_3658_),
    .Z(_0393_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7371_ (.I(\mod.Data_Mem.F_M.MRAM[773][2] ),
    .Z(_3659_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7372_ (.I(_3659_),
    .Z(_0394_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7373_ (.I(\mod.Data_Mem.F_M.MRAM[773][3] ),
    .Z(_3660_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7374_ (.I(_3660_),
    .Z(_0395_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7375_ (.I(\mod.Data_Mem.F_M.MRAM[773][4] ),
    .Z(_3661_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7376_ (.I(_3661_),
    .Z(_0396_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7377_ (.I(\mod.Data_Mem.F_M.MRAM[773][5] ),
    .Z(_3662_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7378_ (.I(_3662_),
    .Z(_0397_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7379_ (.I(\mod.Data_Mem.F_M.MRAM[773][6] ),
    .Z(_3663_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7380_ (.I(_3663_),
    .Z(_0398_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7381_ (.I(\mod.Data_Mem.F_M.MRAM[773][7] ),
    .Z(_3664_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7382_ (.I(_3664_),
    .Z(_0399_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7383_ (.I(\mod.Data_Mem.F_M.MRAM[774][0] ),
    .Z(_3665_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7384_ (.I(_3665_),
    .Z(_0400_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7385_ (.I(\mod.Data_Mem.F_M.MRAM[774][1] ),
    .Z(_3666_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7386_ (.I(_3666_),
    .Z(_0401_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7387_ (.I(\mod.Data_Mem.F_M.MRAM[774][2] ),
    .Z(_3667_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7388_ (.I(_3667_),
    .Z(_0402_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7389_ (.I(\mod.Data_Mem.F_M.MRAM[774][3] ),
    .Z(_3668_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7390_ (.I(_3668_),
    .Z(_0403_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7391_ (.I(\mod.Data_Mem.F_M.MRAM[774][4] ),
    .Z(_3669_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7392_ (.I(_3669_),
    .Z(_0404_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7393_ (.I(\mod.Data_Mem.F_M.MRAM[774][5] ),
    .Z(_3670_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7394_ (.I(_3670_),
    .Z(_0405_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7395_ (.I(\mod.Data_Mem.F_M.MRAM[774][6] ),
    .Z(_3671_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7396_ (.I(_3671_),
    .Z(_0406_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7397_ (.I(\mod.Data_Mem.F_M.MRAM[774][7] ),
    .Z(_3672_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7398_ (.I(_3672_),
    .Z(_0407_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7399_ (.I(\mod.Data_Mem.F_M.MRAM[775][0] ),
    .Z(_3673_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7400_ (.I(_3673_),
    .Z(_0408_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7401_ (.I(\mod.Data_Mem.F_M.MRAM[775][1] ),
    .Z(_3674_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7402_ (.I(_3674_),
    .Z(_0409_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7403_ (.I(\mod.Data_Mem.F_M.MRAM[775][2] ),
    .Z(_3675_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7404_ (.I(_3675_),
    .Z(_0410_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7405_ (.I(\mod.Data_Mem.F_M.MRAM[775][3] ),
    .Z(_3676_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7406_ (.I(_3676_),
    .Z(_0411_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7407_ (.I(\mod.Data_Mem.F_M.MRAM[775][4] ),
    .Z(_3677_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7408_ (.I(_3677_),
    .Z(_0412_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7409_ (.I(\mod.Data_Mem.F_M.MRAM[775][5] ),
    .Z(_3678_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7410_ (.I(_3678_),
    .Z(_0413_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7411_ (.I(\mod.Data_Mem.F_M.MRAM[775][6] ),
    .Z(_3679_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7412_ (.I(_3679_),
    .Z(_0414_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7413_ (.I(\mod.Data_Mem.F_M.MRAM[775][7] ),
    .Z(_3680_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7414_ (.I(_3680_),
    .Z(_0415_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7415_ (.I(\mod.Data_Mem.F_M.MRAM[776][0] ),
    .Z(_3681_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7416_ (.I(_3681_),
    .Z(_0416_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7417_ (.I(\mod.Data_Mem.F_M.MRAM[776][1] ),
    .Z(_3682_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7418_ (.I(_3682_),
    .Z(_0417_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7419_ (.I(\mod.Data_Mem.F_M.MRAM[776][2] ),
    .Z(_3683_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7420_ (.I(_3683_),
    .Z(_0418_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7421_ (.I(\mod.Data_Mem.F_M.MRAM[776][3] ),
    .Z(_3684_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7422_ (.I(_3684_),
    .Z(_0419_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7423_ (.I(\mod.Data_Mem.F_M.MRAM[776][4] ),
    .Z(_3685_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7424_ (.I(_3685_),
    .Z(_0420_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7425_ (.I(\mod.Data_Mem.F_M.MRAM[776][5] ),
    .Z(_3686_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7426_ (.I(_3686_),
    .Z(_0421_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7427_ (.I(\mod.Data_Mem.F_M.MRAM[776][6] ),
    .Z(_3687_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7428_ (.I(_3687_),
    .Z(_0422_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7429_ (.I(\mod.Data_Mem.F_M.MRAM[776][7] ),
    .Z(_3688_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7430_ (.I(_3688_),
    .Z(_0423_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7431_ (.I(\mod.Data_Mem.F_M.MRAM[777][0] ),
    .Z(_3689_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7432_ (.I(_3689_),
    .Z(_0424_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7433_ (.I(\mod.Data_Mem.F_M.MRAM[777][1] ),
    .Z(_3690_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7434_ (.I(_3690_),
    .Z(_0425_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7435_ (.I(\mod.Data_Mem.F_M.MRAM[777][2] ),
    .Z(_3691_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7436_ (.I(_3691_),
    .Z(_0426_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7437_ (.I(\mod.Data_Mem.F_M.MRAM[777][3] ),
    .Z(_3692_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7438_ (.I(_3692_),
    .Z(_0427_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7439_ (.I(\mod.Data_Mem.F_M.MRAM[777][4] ),
    .Z(_3693_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7440_ (.I(_3693_),
    .Z(_0428_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7441_ (.I(\mod.Data_Mem.F_M.MRAM[777][5] ),
    .Z(_3694_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7442_ (.I(_3694_),
    .Z(_0429_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7443_ (.I(\mod.Data_Mem.F_M.MRAM[777][6] ),
    .Z(_3695_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7444_ (.I(_3695_),
    .Z(_0430_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7445_ (.I(\mod.Data_Mem.F_M.MRAM[777][7] ),
    .Z(_3696_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7446_ (.I(_3696_),
    .Z(_0431_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7447_ (.I(\mod.Data_Mem.F_M.MRAM[778][0] ),
    .Z(_3697_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7448_ (.I(_3697_),
    .Z(_0432_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7449_ (.I(\mod.Data_Mem.F_M.MRAM[778][1] ),
    .Z(_3698_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7450_ (.I(_3698_),
    .Z(_0433_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7451_ (.I(\mod.Data_Mem.F_M.MRAM[778][2] ),
    .Z(_3699_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7452_ (.I(_3699_),
    .Z(_0434_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7453_ (.I(\mod.Data_Mem.F_M.MRAM[778][3] ),
    .Z(_3700_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7454_ (.I(_3700_),
    .Z(_0435_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7455_ (.I(\mod.Data_Mem.F_M.MRAM[778][4] ),
    .Z(_3701_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7456_ (.I(_3701_),
    .Z(_0436_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7457_ (.I(\mod.Data_Mem.F_M.MRAM[778][5] ),
    .Z(_3702_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7458_ (.I(_3702_),
    .Z(_0437_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7459_ (.I(\mod.Data_Mem.F_M.MRAM[778][6] ),
    .Z(_3703_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7460_ (.I(_3703_),
    .Z(_0438_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7461_ (.I(\mod.Data_Mem.F_M.MRAM[778][7] ),
    .Z(_3704_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7462_ (.I(_3704_),
    .Z(_0439_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7463_ (.I(_3297_),
    .Z(_3705_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _7464_ (.A1(_3269_),
    .A2(_3705_),
    .A3(_3374_),
    .ZN(_3706_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _7465_ (.I(_3706_),
    .Z(_3707_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _7466_ (.I0(_3603_),
    .I1(\mod.Data_Mem.F_M.MRAM[780][0] ),
    .S(_3707_),
    .Z(_3708_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7467_ (.I(_3708_),
    .Z(_0440_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _7468_ (.I0(_3638_),
    .I1(\mod.Data_Mem.F_M.MRAM[780][1] ),
    .S(_3707_),
    .Z(_3709_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7469_ (.I(_3709_),
    .Z(_0441_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _7470_ (.I0(_3640_),
    .I1(\mod.Data_Mem.F_M.MRAM[780][2] ),
    .S(_3707_),
    .Z(_3710_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7471_ (.I(_3710_),
    .Z(_0442_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7472_ (.I(_3308_),
    .Z(_3711_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _7473_ (.I0(_3711_),
    .I1(\mod.Data_Mem.F_M.MRAM[780][3] ),
    .S(_3707_),
    .Z(_3712_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7474_ (.I(_3712_),
    .Z(_0443_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _7475_ (.I(_3706_),
    .Z(_3713_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _7476_ (.I0(_3615_),
    .I1(\mod.Data_Mem.F_M.MRAM[780][4] ),
    .S(_3713_),
    .Z(_3714_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7477_ (.I(_3714_),
    .Z(_0444_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _7478_ (.I0(_3645_),
    .I1(\mod.Data_Mem.F_M.MRAM[780][5] ),
    .S(_3713_),
    .Z(_3715_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7479_ (.I(_3715_),
    .Z(_0445_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _7480_ (.I0(_3618_),
    .I1(\mod.Data_Mem.F_M.MRAM[780][6] ),
    .S(_3713_),
    .Z(_3716_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7481_ (.I(_3716_),
    .Z(_0446_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _7482_ (.I0(_3620_),
    .I1(\mod.Data_Mem.F_M.MRAM[780][7] ),
    .S(_3713_),
    .Z(_3717_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7483_ (.I(_3717_),
    .Z(_0447_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7484_ (.I(_3292_),
    .Z(_3718_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _7485_ (.A1(_3634_),
    .A2(_3371_),
    .A3(_3387_),
    .ZN(_3719_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _7486_ (.I(_3719_),
    .Z(_3720_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _7487_ (.I0(_3718_),
    .I1(\mod.Data_Mem.F_M.MRAM[781][0] ),
    .S(_3720_),
    .Z(_3721_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7488_ (.I(_3721_),
    .Z(_0448_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _7489_ (.I0(_3638_),
    .I1(\mod.Data_Mem.F_M.MRAM[781][1] ),
    .S(_3720_),
    .Z(_3722_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7490_ (.I(_3722_),
    .Z(_0449_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _7491_ (.I0(_3640_),
    .I1(\mod.Data_Mem.F_M.MRAM[781][2] ),
    .S(_3720_),
    .Z(_3723_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7492_ (.I(_3723_),
    .Z(_0450_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _7493_ (.I0(_3711_),
    .I1(\mod.Data_Mem.F_M.MRAM[781][3] ),
    .S(_3720_),
    .Z(_3724_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7494_ (.I(_3724_),
    .Z(_0451_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7495_ (.I(_3311_),
    .Z(_3725_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _7496_ (.I(_3719_),
    .Z(_3726_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _7497_ (.I0(_3725_),
    .I1(\mod.Data_Mem.F_M.MRAM[781][4] ),
    .S(_3726_),
    .Z(_3727_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7498_ (.I(_3727_),
    .Z(_0452_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _7499_ (.I0(_3645_),
    .I1(\mod.Data_Mem.F_M.MRAM[781][5] ),
    .S(_3726_),
    .Z(_3728_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7500_ (.I(_3728_),
    .Z(_0453_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7501_ (.I(_3318_),
    .Z(_3729_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _7502_ (.I0(_3729_),
    .I1(\mod.Data_Mem.F_M.MRAM[781][6] ),
    .S(_3726_),
    .Z(_3730_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7503_ (.I(_3730_),
    .Z(_0454_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7504_ (.I(_3321_),
    .Z(_3731_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _7505_ (.I0(_3731_),
    .I1(\mod.Data_Mem.F_M.MRAM[781][7] ),
    .S(_3726_),
    .Z(_3732_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7506_ (.I(_3732_),
    .Z(_0455_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _7507_ (.A1(_3634_),
    .A2(_3387_),
    .A3(_3389_),
    .ZN(_3733_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _7508_ (.I(_3733_),
    .Z(_3734_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _7509_ (.I0(_3718_),
    .I1(\mod.Data_Mem.F_M.MRAM[782][0] ),
    .S(_3734_),
    .Z(_3735_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7510_ (.I(_3735_),
    .Z(_0456_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _7511_ (.I0(_3638_),
    .I1(\mod.Data_Mem.F_M.MRAM[782][1] ),
    .S(_3734_),
    .Z(_3736_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7512_ (.I(_3736_),
    .Z(_0457_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _7513_ (.I0(_3640_),
    .I1(\mod.Data_Mem.F_M.MRAM[782][2] ),
    .S(_3734_),
    .Z(_3737_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7514_ (.I(_3737_),
    .Z(_0458_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _7515_ (.I0(_3711_),
    .I1(\mod.Data_Mem.F_M.MRAM[782][3] ),
    .S(_3734_),
    .Z(_3738_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7516_ (.I(_3738_),
    .Z(_0459_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _7517_ (.I(_3733_),
    .Z(_3739_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _7518_ (.I0(_3725_),
    .I1(\mod.Data_Mem.F_M.MRAM[782][4] ),
    .S(_3739_),
    .Z(_3740_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7519_ (.I(_3740_),
    .Z(_0460_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _7520_ (.I0(_3645_),
    .I1(\mod.Data_Mem.F_M.MRAM[782][5] ),
    .S(_3739_),
    .Z(_3741_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7521_ (.I(_3741_),
    .Z(_0461_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _7522_ (.I0(_3729_),
    .I1(\mod.Data_Mem.F_M.MRAM[782][6] ),
    .S(_3739_),
    .Z(_3742_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7523_ (.I(_3742_),
    .Z(_0462_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _7524_ (.I0(_3731_),
    .I1(\mod.Data_Mem.F_M.MRAM[782][7] ),
    .S(_3739_),
    .Z(_3743_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7525_ (.I(_3743_),
    .Z(_0463_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _7526_ (.A1(_3407_),
    .A2(_3705_),
    .A3(_3387_),
    .ZN(_3744_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _7527_ (.I(_3744_),
    .Z(_3745_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _7528_ (.I0(_3718_),
    .I1(\mod.Data_Mem.F_M.MRAM[783][0] ),
    .S(_3745_),
    .Z(_3746_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7529_ (.I(_3746_),
    .Z(_0464_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7530_ (.I(_3302_),
    .Z(_3747_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _7531_ (.I0(_3747_),
    .I1(\mod.Data_Mem.F_M.MRAM[783][1] ),
    .S(_3745_),
    .Z(_3748_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7532_ (.I(_3748_),
    .Z(_0465_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7533_ (.I(_3305_),
    .Z(_3749_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _7534_ (.I0(_3749_),
    .I1(\mod.Data_Mem.F_M.MRAM[783][2] ),
    .S(_3745_),
    .Z(_3750_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7535_ (.I(_3750_),
    .Z(_0466_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _7536_ (.I0(_3711_),
    .I1(\mod.Data_Mem.F_M.MRAM[783][3] ),
    .S(_3745_),
    .Z(_3751_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7537_ (.I(_3751_),
    .Z(_0467_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _7538_ (.I(_3744_),
    .Z(_3752_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _7539_ (.I0(_3725_),
    .I1(_1901_),
    .S(_3752_),
    .Z(_3753_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7540_ (.I(_3753_),
    .Z(_0468_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7541_ (.I(_3315_),
    .Z(_3754_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _7542_ (.I0(_3754_),
    .I1(\mod.Data_Mem.F_M.MRAM[783][5] ),
    .S(_3752_),
    .Z(_3755_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7543_ (.I(_3755_),
    .Z(_0469_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _7544_ (.I0(_3729_),
    .I1(\mod.Data_Mem.F_M.MRAM[783][6] ),
    .S(_3752_),
    .Z(_3756_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7545_ (.I(_3756_),
    .Z(_0470_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _7546_ (.I0(_3731_),
    .I1(\mod.Data_Mem.F_M.MRAM[783][7] ),
    .S(_3752_),
    .Z(_3757_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7547_ (.I(_3757_),
    .Z(_0471_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _7548_ (.I(_3420_),
    .Z(_3758_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _7549_ (.A1(_3232_),
    .A2(_3298_),
    .A3(_3758_),
    .ZN(_3759_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _7550_ (.I(_3759_),
    .Z(_3760_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _7551_ (.I0(_3718_),
    .I1(\mod.Data_Mem.F_M.MRAM[784][0] ),
    .S(_3760_),
    .Z(_3761_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7552_ (.I(_3761_),
    .Z(_0472_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7553_ (.I(_3759_),
    .Z(_3762_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7554_ (.A1(_3610_),
    .A2(_3762_),
    .ZN(_3763_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7555_ (.A1(_1678_),
    .A2(_3762_),
    .B(_3763_),
    .ZN(_0473_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7556_ (.A1(_3612_),
    .A2(_3762_),
    .ZN(_3764_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7557_ (.A1(_1792_),
    .A2(_3762_),
    .B(_3764_),
    .ZN(_0474_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7558_ (.I(_3308_),
    .Z(_3765_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _7559_ (.I0(_3765_),
    .I1(\mod.Data_Mem.F_M.MRAM[784][3] ),
    .S(_3760_),
    .Z(_3766_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7560_ (.I(_3766_),
    .Z(_0475_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _7561_ (.I0(_3725_),
    .I1(\mod.Data_Mem.F_M.MRAM[784][4] ),
    .S(_3760_),
    .Z(_3767_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7562_ (.I(_3767_),
    .Z(_0476_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _7563_ (.I0(_3754_),
    .I1(\mod.Data_Mem.F_M.MRAM[784][5] ),
    .S(_3760_),
    .Z(_3768_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7564_ (.I(_3768_),
    .Z(_0477_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _7565_ (.I0(_3729_),
    .I1(\mod.Data_Mem.F_M.MRAM[784][6] ),
    .S(_3759_),
    .Z(_3769_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7566_ (.I(_3769_),
    .Z(_0478_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _7567_ (.I0(_3731_),
    .I1(\mod.Data_Mem.F_M.MRAM[784][7] ),
    .S(_3759_),
    .Z(_3770_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7568_ (.I(_3770_),
    .Z(_0479_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7569_ (.I(_3292_),
    .Z(_3771_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _7570_ (.A1(_3705_),
    .A2(_3335_),
    .A3(_3758_),
    .ZN(_3772_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _7571_ (.I(_3772_),
    .Z(_3773_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _7572_ (.I0(_3771_),
    .I1(\mod.Data_Mem.F_M.MRAM[785][0] ),
    .S(_3773_),
    .Z(_3774_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7573_ (.I(_3774_),
    .Z(_0480_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _7574_ (.I0(_3747_),
    .I1(\mod.Data_Mem.F_M.MRAM[785][1] ),
    .S(_3773_),
    .Z(_3775_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7575_ (.I(_3775_),
    .Z(_0481_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _7576_ (.I0(_3749_),
    .I1(\mod.Data_Mem.F_M.MRAM[785][2] ),
    .S(_3773_),
    .Z(_3776_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7577_ (.I(_3776_),
    .Z(_0482_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _7578_ (.I0(_3765_),
    .I1(\mod.Data_Mem.F_M.MRAM[785][3] ),
    .S(_3773_),
    .Z(_3777_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7579_ (.I(_3777_),
    .Z(_0483_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7580_ (.I(_3311_),
    .Z(_3778_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _7581_ (.I(_3772_),
    .Z(_3779_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _7582_ (.I0(_3778_),
    .I1(\mod.Data_Mem.F_M.MRAM[785][4] ),
    .S(_3779_),
    .Z(_3780_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7583_ (.I(_3780_),
    .Z(_0484_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _7584_ (.I0(_3754_),
    .I1(\mod.Data_Mem.F_M.MRAM[785][5] ),
    .S(_3779_),
    .Z(_3781_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7585_ (.I(_3781_),
    .Z(_0485_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7586_ (.I(_3318_),
    .Z(_3782_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _7587_ (.I0(_3782_),
    .I1(\mod.Data_Mem.F_M.MRAM[785][6] ),
    .S(_3779_),
    .Z(_3783_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7588_ (.I(_3783_),
    .Z(_0486_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7589_ (.I(_3321_),
    .Z(_3784_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _7590_ (.I0(_3784_),
    .I1(\mod.Data_Mem.F_M.MRAM[785][7] ),
    .S(_3779_),
    .Z(_3785_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7591_ (.I(_3785_),
    .Z(_0487_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_4 _7592_ (.A1(_3604_),
    .A2(_3446_),
    .A3(_3758_),
    .ZN(_3786_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _7593_ (.I(_3786_),
    .Z(_3787_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _7594_ (.I0(_3771_),
    .I1(\mod.Data_Mem.F_M.MRAM[786][0] ),
    .S(_3787_),
    .Z(_3788_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7595_ (.I(_3788_),
    .Z(_0488_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7596_ (.I(_3786_),
    .Z(_3789_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7597_ (.A1(_3610_),
    .A2(_3789_),
    .ZN(_3790_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7598_ (.A1(_1682_),
    .A2(_3789_),
    .B(_3790_),
    .ZN(_0489_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7599_ (.A1(_3612_),
    .A2(_3789_),
    .ZN(_3791_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7600_ (.A1(_1787_),
    .A2(_3789_),
    .B(_3791_),
    .ZN(_0490_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _7601_ (.I0(_3765_),
    .I1(\mod.Data_Mem.F_M.MRAM[786][3] ),
    .S(_3787_),
    .Z(_3792_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7602_ (.I(_3792_),
    .Z(_0491_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _7603_ (.I0(_3778_),
    .I1(\mod.Data_Mem.F_M.MRAM[786][4] ),
    .S(_3787_),
    .Z(_3793_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7604_ (.I(_3793_),
    .Z(_0492_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _7605_ (.I0(_3754_),
    .I1(\mod.Data_Mem.F_M.MRAM[786][5] ),
    .S(_3787_),
    .Z(_3794_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7606_ (.I(_3794_),
    .Z(_0493_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _7607_ (.I0(_3782_),
    .I1(\mod.Data_Mem.F_M.MRAM[786][6] ),
    .S(_3786_),
    .Z(_3795_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7608_ (.I(_3795_),
    .Z(_0494_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _7609_ (.I0(_3784_),
    .I1(\mod.Data_Mem.F_M.MRAM[786][7] ),
    .S(_3786_),
    .Z(_3796_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7610_ (.I(_3796_),
    .Z(_0495_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _7611_ (.A1(_3296_),
    .A2(_3604_),
    .A3(_3758_),
    .ZN(_3797_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7612_ (.I(_3797_),
    .Z(_3798_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _7613_ (.I0(_3771_),
    .I1(\mod.Data_Mem.F_M.MRAM[787][0] ),
    .S(_3798_),
    .Z(_3799_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7614_ (.I(_3799_),
    .Z(_0496_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _7615_ (.I0(_3747_),
    .I1(\mod.Data_Mem.F_M.MRAM[787][1] ),
    .S(_3798_),
    .Z(_3800_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7616_ (.I(_3800_),
    .Z(_0497_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _7617_ (.I(_3797_),
    .Z(_3801_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _7618_ (.I0(_3749_),
    .I1(\mod.Data_Mem.F_M.MRAM[787][2] ),
    .S(_3801_),
    .Z(_3802_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7619_ (.I(_3802_),
    .Z(_0498_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _7620_ (.I0(_3765_),
    .I1(\mod.Data_Mem.F_M.MRAM[787][3] ),
    .S(_3801_),
    .Z(_3803_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7621_ (.I(_3803_),
    .Z(_0499_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7622_ (.I(_3801_),
    .Z(_3804_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7623_ (.A1(_3312_),
    .A2(_3804_),
    .ZN(_3805_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7624_ (.A1(_1919_),
    .A2(_3804_),
    .B(_3805_),
    .ZN(_0500_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7625_ (.I(_3315_),
    .Z(_3806_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _7626_ (.I0(_3806_),
    .I1(\mod.Data_Mem.F_M.MRAM[787][5] ),
    .S(_3801_),
    .Z(_3807_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7627_ (.I(_3807_),
    .Z(_0501_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7628_ (.A1(_3319_),
    .A2(_3798_),
    .ZN(_3808_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7629_ (.A1(_2013_),
    .A2(_3804_),
    .B(_3808_),
    .ZN(_0502_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7630_ (.A1(_3322_),
    .A2(_3798_),
    .ZN(_3809_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7631_ (.A1(_2049_),
    .A2(_3804_),
    .B(_3809_),
    .ZN(_0503_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7632_ (.I(\mod.Data_Mem.F_M.MRAM[788][0] ),
    .Z(_3810_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7633_ (.I(_3810_),
    .Z(_0504_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7634_ (.I(\mod.Data_Mem.F_M.MRAM[788][1] ),
    .Z(_3811_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7635_ (.I(_3811_),
    .Z(_0505_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7636_ (.I(\mod.Data_Mem.F_M.MRAM[788][2] ),
    .Z(_3812_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7637_ (.I(_3812_),
    .Z(_0506_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7638_ (.I(\mod.Data_Mem.F_M.MRAM[788][3] ),
    .Z(_3813_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7639_ (.I(_3813_),
    .Z(_0507_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7640_ (.I(\mod.Data_Mem.F_M.MRAM[788][4] ),
    .Z(_3814_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7641_ (.I(_3814_),
    .Z(_0508_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7642_ (.I(\mod.Data_Mem.F_M.MRAM[788][5] ),
    .Z(_3815_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7643_ (.I(_3815_),
    .Z(_0509_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7644_ (.I(\mod.Data_Mem.F_M.MRAM[788][6] ),
    .Z(_3816_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7645_ (.I(_3816_),
    .Z(_0510_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7646_ (.I(\mod.Data_Mem.F_M.MRAM[788][7] ),
    .Z(_3817_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7647_ (.I(_3817_),
    .Z(_0511_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7648_ (.I(\mod.Data_Mem.F_M.MRAM[790][0] ),
    .Z(_3818_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7649_ (.I(_3818_),
    .Z(_0512_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7650_ (.I(\mod.Data_Mem.F_M.MRAM[790][1] ),
    .Z(_3819_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7651_ (.I(_3819_),
    .Z(_0513_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7652_ (.I(\mod.Data_Mem.F_M.MRAM[790][2] ),
    .Z(_3820_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7653_ (.I(_3820_),
    .Z(_0514_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7654_ (.I(\mod.Data_Mem.F_M.MRAM[790][3] ),
    .Z(_3821_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7655_ (.I(_3821_),
    .Z(_0515_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7656_ (.I(\mod.Data_Mem.F_M.MRAM[790][4] ),
    .Z(_3822_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7657_ (.I(_3822_),
    .Z(_0516_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7658_ (.I(\mod.Data_Mem.F_M.MRAM[790][5] ),
    .Z(_3823_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7659_ (.I(_3823_),
    .Z(_0517_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7660_ (.I(\mod.Data_Mem.F_M.MRAM[790][6] ),
    .Z(_3824_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7661_ (.I(_3824_),
    .Z(_0518_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7662_ (.I(\mod.Data_Mem.F_M.MRAM[790][7] ),
    .Z(_3825_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7663_ (.I(_3825_),
    .Z(_0519_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7664_ (.I(\mod.Data_Mem.F_M.MRAM[791][0] ),
    .Z(_3826_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7665_ (.I(_3826_),
    .Z(_0520_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7666_ (.I(\mod.Data_Mem.F_M.MRAM[791][1] ),
    .Z(_3827_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7667_ (.I(_3827_),
    .Z(_0521_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7668_ (.I(\mod.Data_Mem.F_M.MRAM[791][2] ),
    .Z(_3828_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7669_ (.I(_3828_),
    .Z(_0522_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7670_ (.I(\mod.Data_Mem.F_M.MRAM[791][3] ),
    .Z(_3829_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7671_ (.I(_3829_),
    .Z(_0523_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7672_ (.I(\mod.Data_Mem.F_M.MRAM[791][4] ),
    .Z(_3830_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7673_ (.I(_3830_),
    .Z(_0524_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7674_ (.I(\mod.Data_Mem.F_M.MRAM[791][5] ),
    .Z(_3831_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7675_ (.I(_3831_),
    .Z(_0525_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7676_ (.I(\mod.Data_Mem.F_M.MRAM[791][6] ),
    .Z(_3832_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7677_ (.I(_3832_),
    .Z(_0526_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7678_ (.I(\mod.Data_Mem.F_M.MRAM[791][7] ),
    .Z(_3833_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7679_ (.I(_3833_),
    .Z(_0527_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7680_ (.I(\mod.Data_Mem.F_M.MRAM[792][0] ),
    .Z(_3834_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7681_ (.I(_3834_),
    .Z(_0528_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7682_ (.I(\mod.Data_Mem.F_M.MRAM[792][1] ),
    .Z(_3835_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7683_ (.I(_3835_),
    .Z(_0529_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7684_ (.I(\mod.Data_Mem.F_M.MRAM[792][2] ),
    .Z(_3836_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7685_ (.I(_3836_),
    .Z(_0530_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7686_ (.I(\mod.Data_Mem.F_M.MRAM[792][3] ),
    .Z(_3837_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7687_ (.I(_3837_),
    .Z(_0531_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7688_ (.I(\mod.Data_Mem.F_M.MRAM[792][4] ),
    .Z(_3838_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7689_ (.I(_3838_),
    .Z(_0532_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7690_ (.I(\mod.Data_Mem.F_M.MRAM[792][5] ),
    .Z(_3839_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7691_ (.I(_3839_),
    .Z(_0533_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7692_ (.I(\mod.Data_Mem.F_M.MRAM[792][6] ),
    .Z(_3840_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7693_ (.I(_3840_),
    .Z(_0534_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7694_ (.I(\mod.Data_Mem.F_M.MRAM[792][7] ),
    .Z(_3841_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7695_ (.I(_3841_),
    .Z(_0535_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7696_ (.I(\mod.Data_Mem.F_M.MRAM[793][0] ),
    .Z(_3842_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7697_ (.I(_3842_),
    .Z(_0536_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7698_ (.I(\mod.Data_Mem.F_M.MRAM[793][1] ),
    .Z(_3843_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7699_ (.I(_3843_),
    .Z(_0537_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7700_ (.I(\mod.Data_Mem.F_M.MRAM[793][2] ),
    .Z(_3844_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7701_ (.I(_3844_),
    .Z(_0538_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7702_ (.I(\mod.Data_Mem.F_M.MRAM[793][3] ),
    .Z(_3845_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7703_ (.I(_3845_),
    .Z(_0539_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7704_ (.I(\mod.Data_Mem.F_M.MRAM[793][4] ),
    .Z(_3846_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7705_ (.I(_3846_),
    .Z(_0540_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7706_ (.I(\mod.Data_Mem.F_M.MRAM[793][5] ),
    .Z(_3847_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7707_ (.I(_3847_),
    .Z(_0541_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7708_ (.I(\mod.Data_Mem.F_M.MRAM[793][6] ),
    .Z(_3848_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7709_ (.I(_3848_),
    .Z(_0542_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7710_ (.I(\mod.Data_Mem.F_M.MRAM[793][7] ),
    .Z(_3849_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7711_ (.I(_3849_),
    .Z(_0543_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7712_ (.I(\mod.Data_Mem.F_M.MRAM[794][0] ),
    .Z(_3850_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7713_ (.I(_3850_),
    .Z(_0544_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7714_ (.I(\mod.Data_Mem.F_M.MRAM[794][1] ),
    .Z(_3851_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7715_ (.I(_3851_),
    .Z(_0545_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7716_ (.I(\mod.Data_Mem.F_M.MRAM[794][2] ),
    .Z(_3852_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7717_ (.I(_3852_),
    .Z(_0546_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7718_ (.I(\mod.Data_Mem.F_M.MRAM[794][3] ),
    .Z(_3853_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7719_ (.I(_3853_),
    .Z(_0547_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7720_ (.I(\mod.Data_Mem.F_M.MRAM[794][4] ),
    .Z(_3854_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7721_ (.I(_3854_),
    .Z(_0548_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7722_ (.I(\mod.Data_Mem.F_M.MRAM[794][5] ),
    .Z(_3855_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7723_ (.I(_3855_),
    .Z(_0549_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7724_ (.I(\mod.Data_Mem.F_M.MRAM[794][6] ),
    .Z(_3856_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7725_ (.I(_3856_),
    .Z(_0550_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7726_ (.I(\mod.Data_Mem.F_M.MRAM[794][7] ),
    .Z(_3857_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7727_ (.I(_3857_),
    .Z(_0551_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7728_ (.I(\mod.Data_Mem.F_M.MRAM[795][0] ),
    .Z(_3858_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7729_ (.I(_3858_),
    .Z(_0552_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7730_ (.I(\mod.Data_Mem.F_M.MRAM[795][1] ),
    .Z(_3859_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7731_ (.I(_3859_),
    .Z(_0553_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7732_ (.I(\mod.Data_Mem.F_M.MRAM[795][2] ),
    .Z(_3860_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7733_ (.I(_3860_),
    .Z(_0554_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7734_ (.I(\mod.Data_Mem.F_M.MRAM[795][3] ),
    .Z(_3861_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7735_ (.I(_3861_),
    .Z(_0555_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7736_ (.I(\mod.Data_Mem.F_M.MRAM[795][4] ),
    .Z(_3862_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7737_ (.I(_3862_),
    .Z(_0556_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7738_ (.I(\mod.Data_Mem.F_M.MRAM[795][5] ),
    .Z(_3863_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7739_ (.I(_3863_),
    .Z(_0557_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7740_ (.I(\mod.Data_Mem.F_M.MRAM[795][6] ),
    .Z(_3864_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7741_ (.I(_3864_),
    .Z(_0558_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7742_ (.I(\mod.Data_Mem.F_M.MRAM[795][7] ),
    .Z(_3865_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7743_ (.I(_3865_),
    .Z(_0559_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _7744_ (.A1(_3230_),
    .A2(_3232_),
    .A3(_3634_),
    .ZN(_3866_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _7745_ (.I(_3866_),
    .Z(_3867_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _7746_ (.I0(_3771_),
    .I1(\mod.Data_Mem.F_M.MRAM[796][0] ),
    .S(_3867_),
    .Z(_3868_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7747_ (.I(_3868_),
    .Z(_0560_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _7748_ (.I0(_3747_),
    .I1(\mod.Data_Mem.F_M.MRAM[796][1] ),
    .S(_3867_),
    .Z(_3869_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7749_ (.I(_3869_),
    .Z(_0561_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _7750_ (.I0(_3749_),
    .I1(\mod.Data_Mem.F_M.MRAM[796][2] ),
    .S(_3867_),
    .Z(_3870_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7751_ (.I(_3870_),
    .Z(_0562_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _7752_ (.I0(_3309_),
    .I1(\mod.Data_Mem.F_M.MRAM[796][3] ),
    .S(_3867_),
    .Z(_3871_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7753_ (.I(_3871_),
    .Z(_0563_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _7754_ (.I(_3866_),
    .Z(_3872_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _7755_ (.I0(_3778_),
    .I1(\mod.Data_Mem.F_M.MRAM[796][4] ),
    .S(_3872_),
    .Z(_3873_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7756_ (.I(_3873_),
    .Z(_0564_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _7757_ (.I0(_3806_),
    .I1(\mod.Data_Mem.F_M.MRAM[796][5] ),
    .S(_3872_),
    .Z(_3874_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7758_ (.I(_3874_),
    .Z(_0565_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _7759_ (.I0(_3782_),
    .I1(\mod.Data_Mem.F_M.MRAM[796][6] ),
    .S(_3872_),
    .Z(_3875_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7760_ (.I(_3875_),
    .Z(_0566_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _7761_ (.I0(_3784_),
    .I1(\mod.Data_Mem.F_M.MRAM[796][7] ),
    .S(_3872_),
    .Z(_3876_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7762_ (.I(_3876_),
    .Z(_0567_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _7763_ (.A1(_3230_),
    .A2(_3705_),
    .A3(_3371_),
    .ZN(_3877_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _7764_ (.I(_3877_),
    .Z(_3878_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _7765_ (.I0(_3293_),
    .I1(\mod.Data_Mem.F_M.MRAM[797][0] ),
    .S(_3878_),
    .Z(_3879_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7766_ (.I(_3879_),
    .Z(_0568_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _7767_ (.I0(_3303_),
    .I1(\mod.Data_Mem.F_M.MRAM[797][1] ),
    .S(_3878_),
    .Z(_3880_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7768_ (.I(_3880_),
    .Z(_0569_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _7769_ (.I0(_3306_),
    .I1(\mod.Data_Mem.F_M.MRAM[797][2] ),
    .S(_3878_),
    .Z(_3881_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7770_ (.I(_3881_),
    .Z(_0570_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _7771_ (.I0(_3309_),
    .I1(\mod.Data_Mem.F_M.MRAM[797][3] ),
    .S(_3878_),
    .Z(_3882_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7772_ (.I(_3882_),
    .Z(_0571_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _7773_ (.I(_3877_),
    .Z(_3883_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _7774_ (.I0(_3778_),
    .I1(\mod.Data_Mem.F_M.MRAM[797][4] ),
    .S(_3883_),
    .Z(_3884_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7775_ (.I(_3884_),
    .Z(_0572_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _7776_ (.I0(_3806_),
    .I1(\mod.Data_Mem.F_M.MRAM[797][5] ),
    .S(_3883_),
    .Z(_3885_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7777_ (.I(_3885_),
    .Z(_0573_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _7778_ (.I0(_3782_),
    .I1(\mod.Data_Mem.F_M.MRAM[797][6] ),
    .S(_3883_),
    .Z(_3886_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7779_ (.I(_3886_),
    .Z(_0574_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _7780_ (.I0(_3784_),
    .I1(\mod.Data_Mem.F_M.MRAM[797][7] ),
    .S(_3883_),
    .Z(_3887_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7781_ (.I(_3887_),
    .Z(_0575_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _7782_ (.A1(_3294_),
    .A2(_3298_),
    .A3(_3446_),
    .ZN(_3888_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _7783_ (.I(_3888_),
    .Z(_3889_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _7784_ (.I0(_3293_),
    .I1(\mod.Data_Mem.F_M.MRAM[798][0] ),
    .S(_3889_),
    .Z(_3890_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7785_ (.I(_3890_),
    .Z(_0576_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _7786_ (.I0(_3303_),
    .I1(\mod.Data_Mem.F_M.MRAM[798][1] ),
    .S(_3889_),
    .Z(_3891_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7787_ (.I(_3891_),
    .Z(_0577_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _7788_ (.I0(_3306_),
    .I1(\mod.Data_Mem.F_M.MRAM[798][2] ),
    .S(_3889_),
    .Z(_3892_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7789_ (.I(_3892_),
    .Z(_0578_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _7790_ (.I0(_3309_),
    .I1(\mod.Data_Mem.F_M.MRAM[798][3] ),
    .S(_3889_),
    .Z(_3893_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7791_ (.I(_3893_),
    .Z(_0579_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _7792_ (.I(_3888_),
    .Z(_3894_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _7793_ (.I0(_3312_),
    .I1(\mod.Data_Mem.F_M.MRAM[798][4] ),
    .S(_3894_),
    .Z(_3895_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7794_ (.I(_3895_),
    .Z(_0580_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _7795_ (.I0(_3806_),
    .I1(\mod.Data_Mem.F_M.MRAM[798][5] ),
    .S(_3894_),
    .Z(_3896_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7796_ (.I(_3896_),
    .Z(_0581_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _7797_ (.I0(_3319_),
    .I1(\mod.Data_Mem.F_M.MRAM[798][6] ),
    .S(_3894_),
    .Z(_3897_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7798_ (.I(_3897_),
    .Z(_0582_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _7799_ (.I0(_3322_),
    .I1(\mod.Data_Mem.F_M.MRAM[798][7] ),
    .S(_3894_),
    .Z(_3898_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7800_ (.I(_3898_),
    .Z(_0583_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7801_ (.I(\mod.Data_Mem.F_M.MRAM[7][0] ),
    .Z(_3899_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7802_ (.I(_3899_),
    .Z(_0584_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7803_ (.I(\mod.Data_Mem.F_M.MRAM[7][1] ),
    .Z(_3900_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7804_ (.I(_3900_),
    .Z(_0585_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7805_ (.I(\mod.Data_Mem.F_M.MRAM[7][2] ),
    .Z(_3901_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7806_ (.I(_3901_),
    .Z(_0586_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7807_ (.I(\mod.Data_Mem.F_M.MRAM[7][3] ),
    .Z(_3902_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7808_ (.I(_3902_),
    .Z(_0587_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7809_ (.I(\mod.Data_Mem.F_M.MRAM[7][4] ),
    .Z(_3903_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7810_ (.I(_3903_),
    .Z(_0588_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7811_ (.I(\mod.Data_Mem.F_M.MRAM[7][5] ),
    .Z(_3904_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7812_ (.I(_3904_),
    .Z(_0589_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7813_ (.I(\mod.Data_Mem.F_M.MRAM[7][6] ),
    .Z(_3905_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7814_ (.I(_3905_),
    .Z(_0590_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7815_ (.I(\mod.Data_Mem.F_M.MRAM[7][7] ),
    .Z(_3906_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7816_ (.I(_3906_),
    .Z(_0591_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7817_ (.I(\mod.I_addr[3] ),
    .Z(_3907_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _7818_ (.A1(\mod.I_addr[4] ),
    .A2(\mod.I_addr[6] ),
    .A3(\mod.I_addr[5] ),
    .A4(\mod.I_addr[7] ),
    .ZN(_3908_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _7819_ (.A1(\mod.I_addr[0] ),
    .A2(\mod.I_addr[2] ),
    .A3(\mod.I_addr[1] ),
    .ZN(_3909_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _7820_ (.A1(_3907_),
    .A2(_3908_),
    .A3(_3909_),
    .Z(_3910_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7821_ (.I(_3910_),
    .Z(_0592_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7822_ (.A1(\mod.I_addr[0] ),
    .A2(_3169_),
    .ZN(_3911_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7823_ (.A1(_3171_),
    .A2(_3908_),
    .ZN(_3912_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _7824_ (.A1(_3907_),
    .A2(_3911_),
    .A3(_3912_),
    .ZN(_0593_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7825_ (.A1(_3907_),
    .A2(_3912_),
    .ZN(_0594_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7826_ (.A1(\mod.I_addr[3] ),
    .A2(_3911_),
    .ZN(_3913_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _7827_ (.A1(_3908_),
    .A2(_3913_),
    .Z(_3914_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7828_ (.I(_3914_),
    .Z(_0595_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7829_ (.A1(_3174_),
    .A2(_3909_),
    .B(_3908_),
    .ZN(_3915_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7830_ (.I(_3915_),
    .Z(_3916_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7831_ (.A1(_0612_),
    .A2(_3175_),
    .B(_3916_),
    .ZN(_0596_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7832_ (.I(_3916_),
    .Z(_3917_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7833_ (.A1(_0081_),
    .A2(_3917_),
    .ZN(_0597_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7834_ (.A1(_0080_),
    .A2(_3171_),
    .Z(_3918_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7835_ (.A1(_3175_),
    .A2(_3918_),
    .B(_3916_),
    .ZN(_0598_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7836_ (.A1(_3907_),
    .A2(\mod.I_addr[2] ),
    .ZN(_3919_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _7837_ (.A1(_3913_),
    .A2(_3915_),
    .A3(_3919_),
    .ZN(_3920_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7838_ (.I(_3920_),
    .Z(_0610_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _7839_ (.I(_3169_),
    .ZN(_3921_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _7840_ (.A1(_0080_),
    .A2(_3171_),
    .B(_3921_),
    .C(_3916_),
    .ZN(_3922_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _7841_ (.A1(_0610_),
    .A2(_3922_),
    .Z(_3923_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7842_ (.I(_3923_),
    .Z(_0599_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7843_ (.I(\mod.Data_Mem.F_M.MRAM[9][0] ),
    .Z(_3924_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7844_ (.I(_3924_),
    .Z(_0600_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7845_ (.I(\mod.Data_Mem.F_M.MRAM[9][1] ),
    .Z(_3925_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7846_ (.I(_3925_),
    .Z(_0601_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7847_ (.I(\mod.Data_Mem.F_M.MRAM[9][2] ),
    .Z(_3926_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7848_ (.I(_3926_),
    .Z(_0602_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7849_ (.I(\mod.Data_Mem.F_M.MRAM[9][3] ),
    .Z(_3927_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7850_ (.I(_3927_),
    .Z(_0603_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7851_ (.I(\mod.Data_Mem.F_M.MRAM[9][4] ),
    .Z(_3928_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7852_ (.I(_3928_),
    .Z(_0604_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7853_ (.I(\mod.Data_Mem.F_M.MRAM[9][5] ),
    .Z(_3929_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7854_ (.I(_3929_),
    .Z(_0605_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7855_ (.I(\mod.Data_Mem.F_M.MRAM[9][6] ),
    .Z(_3930_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7856_ (.I(_3930_),
    .Z(_0606_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7857_ (.I(\mod.Data_Mem.F_M.MRAM[9][7] ),
    .Z(_3931_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7858_ (.I(_3931_),
    .Z(_0607_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7859_ (.A1(_3913_),
    .A2(_3917_),
    .ZN(_0608_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _7860_ (.I(_3917_),
    .ZN(_0609_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7861_ (.A1(_3917_),
    .A2(_3919_),
    .ZN(_0611_));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7862_ (.D(_0088_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.MRAM[11][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7863_ (.D(_0089_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.MRAM[11][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7864_ (.D(_0090_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.MRAM[11][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7865_ (.D(_0091_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.MRAM[11][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7866_ (.D(_0092_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.MRAM[11][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7867_ (.D(_0093_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.MRAM[11][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7868_ (.D(_0094_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.MRAM[11][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7869_ (.D(_0095_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.MRAM[11][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7870_ (.D(_0096_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.MRAM[24][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7871_ (.D(_0097_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.MRAM[24][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7872_ (.D(_0098_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.MRAM[24][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7873_ (.D(_0099_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.MRAM[24][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7874_ (.D(_0100_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.MRAM[24][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7875_ (.D(_0101_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.MRAM[24][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7876_ (.D(_0102_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.MRAM[24][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7877_ (.D(_0103_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.MRAM[24][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7878_ (.D(_0104_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.MRAM[26][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7879_ (.D(_0105_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.MRAM[26][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7880_ (.D(_0106_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.MRAM[26][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7881_ (.D(_0107_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.MRAM[26][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7882_ (.D(_0108_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.MRAM[26][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7883_ (.D(_0109_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.MRAM[26][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7884_ (.D(_0110_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.MRAM[26][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7885_ (.D(_0111_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.MRAM[26][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7886_ (.D(_0112_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.MRAM[25][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7887_ (.D(_0113_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.MRAM[25][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7888_ (.D(_0114_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.MRAM[25][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7889_ (.D(_0115_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.MRAM[25][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7890_ (.D(_0116_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.MRAM[25][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7891_ (.D(_0117_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.MRAM[25][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7892_ (.D(_0118_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.MRAM[25][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7893_ (.D(_0119_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.MRAM[25][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7894_ (.D(_0120_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.MRAM[27][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7895_ (.D(_0121_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.MRAM[27][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7896_ (.D(_0122_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.MRAM[27][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7897_ (.D(_0123_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.MRAM[27][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7898_ (.D(_0124_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.MRAM[27][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7899_ (.D(_0125_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.MRAM[27][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7900_ (.D(_0126_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.MRAM[27][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7901_ (.D(_0127_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.MRAM[27][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7902_ (.D(_0128_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.MRAM[28][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7903_ (.D(_0129_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.MRAM[28][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7904_ (.D(_0130_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.MRAM[28][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7905_ (.D(_0131_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.MRAM[28][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7906_ (.D(_0132_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.MRAM[28][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7907_ (.D(_0133_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.MRAM[28][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7908_ (.D(_0134_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.MRAM[28][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7909_ (.D(_0135_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.MRAM[28][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7910_ (.D(_0136_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.MRAM[10][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7911_ (.D(_0137_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.MRAM[10][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7912_ (.D(_0138_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.MRAM[10][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7913_ (.D(_0139_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.MRAM[10][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7914_ (.D(_0140_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.MRAM[10][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7915_ (.D(_0141_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.MRAM[10][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7916_ (.D(_0142_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.MRAM[10][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7917_ (.D(_0143_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.MRAM[10][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7918_ (.D(_0144_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.MRAM[0][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7919_ (.D(_0145_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.MRAM[0][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7920_ (.D(_0146_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.MRAM[0][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7921_ (.D(_0147_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.MRAM[0][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7922_ (.D(_0148_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.MRAM[0][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7923_ (.D(_0149_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.MRAM[0][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7924_ (.D(_0150_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.MRAM[0][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7925_ (.D(_0151_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.MRAM[0][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7926_ (.D(_0152_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.MRAM[8][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7927_ (.D(_0153_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.MRAM[8][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7928_ (.D(_0154_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.MRAM[8][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7929_ (.D(_0155_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.MRAM[8][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7930_ (.D(_0156_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.MRAM[8][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7931_ (.D(_0157_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.MRAM[8][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7932_ (.D(_0158_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.MRAM[8][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7933_ (.D(_0159_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.MRAM[8][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7934_ (.D(_0160_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.MRAM[799][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7935_ (.D(_0161_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.MRAM[799][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7936_ (.D(_0162_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.MRAM[799][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7937_ (.D(_0163_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.MRAM[799][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7938_ (.D(_0164_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.MRAM[799][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7939_ (.D(_0165_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.MRAM[799][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7940_ (.D(_0166_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.MRAM[799][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7941_ (.D(_0167_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.MRAM[799][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7942_ (.D(_0168_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.MRAM[789][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7943_ (.D(_0169_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.MRAM[789][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7944_ (.D(_0170_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.MRAM[789][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7945_ (.D(_0171_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.MRAM[789][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7946_ (.D(_0172_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.MRAM[789][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7947_ (.D(_0173_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.MRAM[789][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7948_ (.D(_0174_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.MRAM[789][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7949_ (.D(_0175_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.MRAM[789][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7950_ (.D(_0176_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.MRAM[769][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7951_ (.D(_0177_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.MRAM[769][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7952_ (.D(_0178_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.MRAM[769][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7953_ (.D(_0179_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.MRAM[769][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7954_ (.D(_0180_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.MRAM[769][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7955_ (.D(_0181_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.MRAM[769][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7956_ (.D(_0182_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.MRAM[769][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7957_ (.D(_0183_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.MRAM[769][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7958_ (.D(_0184_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.MRAM[779][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7959_ (.D(_0185_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.MRAM[779][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7960_ (.D(_0186_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.MRAM[779][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7961_ (.D(_0187_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.MRAM[779][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7962_ (.D(_0188_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.MRAM[779][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7963_ (.D(_0189_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.MRAM[779][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7964_ (.D(_0190_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.MRAM[779][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7965_ (.D(_0191_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.MRAM[779][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7966_ (.D(_0192_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.MRAM[6][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7967_ (.D(_0193_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.MRAM[6][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7968_ (.D(_0194_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.MRAM[6][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7969_ (.D(_0195_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.MRAM[6][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7970_ (.D(_0196_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.MRAM[6][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7971_ (.D(_0197_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.MRAM[6][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7972_ (.D(_0198_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.MRAM[6][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7973_ (.D(_0199_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.MRAM[6][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7974_ (.D(_0200_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.MRAM[4][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7975_ (.D(_0201_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.MRAM[4][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7976_ (.D(_0202_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.MRAM[4][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7977_ (.D(_0203_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.MRAM[4][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7978_ (.D(_0204_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.MRAM[4][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7979_ (.D(_0205_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.MRAM[4][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7980_ (.D(_0206_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.MRAM[4][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7981_ (.D(_0207_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.MRAM[4][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _7982_ (.D(\mod.Instr_Mem.instruction[7] ),
    .RN(net2),
    .CLK(net1),
    .Q(\mod.P1.instr_reg[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _7983_ (.D(\mod.Instr_Mem.instruction[8] ),
    .RN(net2),
    .CLK(net1),
    .Q(\mod.P1.instr_reg[8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _7984_ (.D(\mod.Instr_Mem.instruction[9] ),
    .RN(net2),
    .CLK(net1),
    .Q(\mod.P1.instr_reg[9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _7985_ (.D(\mod.Instr_Mem.instruction[10] ),
    .RN(net2),
    .CLK(net1),
    .Q(\mod.P1.instr_reg[10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _7986_ (.D(\mod.Instr_Mem.instruction[11] ),
    .RN(net2),
    .CLK(net1),
    .Q(\mod.P1.instr_reg[11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _7987_ (.D(\mod.Instr_Mem.instruction[13] ),
    .RN(net2),
    .CLK(net1),
    .Q(\mod.P1.instr_reg[13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _7988_ (.D(\mod.Instr_Mem.instruction[17] ),
    .RN(net2),
    .CLK(net1),
    .Q(\mod.P1.instr_reg[17] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _7989_ (.D(\mod.Instr_Mem.instruction[22] ),
    .RN(net2),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.src[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _7990_ (.D(\mod.Instr_Mem.instruction[23] ),
    .RN(net2),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.src[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _7991_ (.D(\mod.Instr_Mem.instruction[24] ),
    .RN(net2),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.src[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _7992_ (.D(\mod.Instr_Mem.instruction[26] ),
    .RN(net2),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.src[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _7993_ (.D(\mod.Instr_Mem.instruction[30] ),
    .RN(net2),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.src[8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _7994_ (.D(\mod.P2.dest_reg1[0] ),
    .RN(net2),
    .CLK(net1),
    .Q(\mod.P2.dest_reg[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _7995_ (.D(\mod.P2.dest_reg1[1] ),
    .RN(net2),
    .CLK(net1),
    .Q(\mod.P2.dest_reg[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _7996_ (.D(\mod.P2.dest_reg1[2] ),
    .RN(net2),
    .CLK(net1),
    .Q(\mod.P2.dest_reg[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _7997_ (.D(\mod.P2.dest_reg1[4] ),
    .RN(net2),
    .CLK(net1),
    .Q(\mod.P2.dest_reg[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _7998_ (.D(\mod.P2.dest_reg1[8] ),
    .RN(net2),
    .CLK(net1),
    .Q(\mod.P2.dest_reg[8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7999_ (.D(_0208_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.MRAM[13][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8000_ (.D(_0209_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.MRAM[13][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8001_ (.D(_0210_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.MRAM[13][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8002_ (.D(_0211_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.MRAM[13][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8003_ (.D(_0212_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.MRAM[13][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8004_ (.D(_0213_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.MRAM[13][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8005_ (.D(_0214_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.MRAM[13][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8006_ (.D(_0215_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.MRAM[13][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8007_ (.D(_0216_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.MRAM[14][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8008_ (.D(_0217_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.MRAM[14][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8009_ (.D(_0218_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.MRAM[14][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8010_ (.D(_0219_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.MRAM[14][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8011_ (.D(_0220_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.MRAM[14][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8012_ (.D(_0221_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.MRAM[14][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8013_ (.D(_0222_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.MRAM[14][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8014_ (.D(_0223_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.MRAM[14][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8015_ (.D(_0224_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.MRAM[15][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8016_ (.D(_0225_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.MRAM[15][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8017_ (.D(_0226_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.MRAM[15][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8018_ (.D(_0227_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.MRAM[15][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8019_ (.D(_0228_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.MRAM[15][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8020_ (.D(_0229_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.MRAM[15][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8021_ (.D(_0230_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.MRAM[15][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8022_ (.D(_0231_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.MRAM[15][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8023_ (.D(_0232_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.MRAM[16][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8024_ (.D(_0233_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.MRAM[16][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8025_ (.D(_0234_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.MRAM[16][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8026_ (.D(_0235_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.MRAM[16][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8027_ (.D(_0236_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.MRAM[16][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8028_ (.D(_0237_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.MRAM[16][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8029_ (.D(_0238_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.MRAM[16][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8030_ (.D(_0239_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.MRAM[16][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8031_ (.D(_0240_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.MRAM[17][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8032_ (.D(_0241_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.MRAM[17][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8033_ (.D(_0242_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.MRAM[17][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8034_ (.D(_0243_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.MRAM[17][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8035_ (.D(_0244_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.MRAM[17][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8036_ (.D(_0245_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.MRAM[17][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8037_ (.D(_0246_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.MRAM[17][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8038_ (.D(_0247_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.MRAM[17][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8039_ (.D(_0248_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.MRAM[18][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8040_ (.D(_0249_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.MRAM[18][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8041_ (.D(_0250_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.MRAM[18][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8042_ (.D(_0251_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.MRAM[18][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8043_ (.D(_0252_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.MRAM[18][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8044_ (.D(_0253_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.MRAM[18][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8045_ (.D(_0254_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.MRAM[18][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8046_ (.D(_0255_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.MRAM[18][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8047_ (.D(_0256_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.MRAM[1][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8048_ (.D(_0257_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.MRAM[1][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8049_ (.D(_0258_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.MRAM[1][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8050_ (.D(_0259_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.MRAM[1][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8051_ (.D(_0260_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.MRAM[1][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8052_ (.D(_0261_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.MRAM[1][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8053_ (.D(_0262_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.MRAM[1][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8054_ (.D(_0263_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.MRAM[1][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8055_ (.D(_0264_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.MRAM[20][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8056_ (.D(_0265_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.MRAM[20][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8057_ (.D(_0266_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.MRAM[20][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8058_ (.D(_0267_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.MRAM[20][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8059_ (.D(_0268_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.MRAM[20][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8060_ (.D(_0269_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.MRAM[20][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8061_ (.D(_0270_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.MRAM[20][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8062_ (.D(_0271_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.MRAM[20][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8063_ (.D(_0272_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.MRAM[21][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8064_ (.D(_0273_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.MRAM[21][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8065_ (.D(_0274_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.MRAM[21][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8066_ (.D(_0275_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.MRAM[21][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8067_ (.D(_0276_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.MRAM[21][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8068_ (.D(_0277_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.MRAM[21][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8069_ (.D(_0278_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.MRAM[21][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8070_ (.D(_0279_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.MRAM[21][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _8071_ (.D(\mod.DMen_reg ),
    .RN(net2),
    .CLK(net1),
    .Q(\mod.DMen_reg2 ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _8072_ (.D(\mod.P3.Res[0] ),
    .RN(net2),
    .CLK(net1),
    .Q(net3));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _8073_ (.D(\mod.P3.Res[1] ),
    .RN(net2),
    .CLK(net1),
    .Q(net4));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _8074_ (.D(\mod.P3.Res[2] ),
    .RN(net2),
    .CLK(net1),
    .Q(net5));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _8075_ (.D(\mod.P3.Res[3] ),
    .RN(net2),
    .CLK(net1),
    .Q(net6));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _8076_ (.D(\mod.P3.Res[4] ),
    .RN(net2),
    .CLK(net1),
    .Q(net7));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _8077_ (.D(\mod.P3.Res[5] ),
    .RN(net2),
    .CLK(net1),
    .Q(net8));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _8078_ (.D(\mod.P3.Res[6] ),
    .RN(net2),
    .CLK(net1),
    .Q(net9));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _8079_ (.D(\mod.P3.Res[7] ),
    .RN(net2),
    .CLK(net1),
    .Q(net10));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8080_ (.D(_0280_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.MRAM[23][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8081_ (.D(_0281_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.MRAM[23][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8082_ (.D(_0282_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.MRAM[23][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8083_ (.D(_0283_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.MRAM[23][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8084_ (.D(_0284_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.MRAM[23][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8085_ (.D(_0285_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.MRAM[23][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8086_ (.D(_0286_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.MRAM[23][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8087_ (.D(_0287_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.MRAM[23][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _8088_ (.D(\mod.P2.Rout_reg1[0] ),
    .RN(net2),
    .CLK(net1),
    .Q(\mod.P2.Rout_reg[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _8089_ (.D(\mod.P2.Rout_reg1[1] ),
    .RN(net2),
    .CLK(net1),
    .Q(\mod.P2.Rout_reg[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _8090_ (.D(\mod.Data_Mem.F_M.out_data[0] ),
    .RN(net2),
    .CLK(net1),
    .Q(\mod.Arithmetic.ACTI.x[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _8091_ (.D(\mod.Data_Mem.F_M.out_data[1] ),
    .RN(net2),
    .CLK(net1),
    .Q(\mod.Arithmetic.ACTI.x[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _8092_ (.D(\mod.Data_Mem.F_M.out_data[2] ),
    .RN(net2),
    .CLK(net1),
    .Q(\mod.Arithmetic.ACTI.x[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _8093_ (.D(\mod.Data_Mem.F_M.out_data[3] ),
    .RN(net2),
    .CLK(net1),
    .Q(\mod.Arithmetic.ACTI.x[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _8094_ (.D(\mod.Data_Mem.F_M.out_data[4] ),
    .RN(net2),
    .CLK(net1),
    .Q(\mod.Arithmetic.ACTI.x[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _8095_ (.D(\mod.Data_Mem.F_M.out_data[5] ),
    .RN(net2),
    .CLK(net1),
    .Q(\mod.Arithmetic.ACTI.x[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _8096_ (.D(\mod.Data_Mem.F_M.out_data[6] ),
    .RN(net2),
    .CLK(net1),
    .Q(\mod.Arithmetic.ACTI.x[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _8097_ (.D(\mod.Data_Mem.F_M.out_data[7] ),
    .RN(net2),
    .CLK(net1),
    .Q(\mod.Arithmetic.ACTI.x[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _8098_ (.D(\mod.Data_Mem.F_M.out_data[8] ),
    .RN(net2),
    .CLK(net1),
    .Q(\mod.Arithmetic.CN.I_in[8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _8099_ (.D(\mod.Data_Mem.F_M.out_data[9] ),
    .RN(net2),
    .CLK(net1),
    .Q(\mod.Arithmetic.CN.I_in[9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _8100_ (.D(\mod.Data_Mem.F_M.out_data[10] ),
    .RN(net2),
    .CLK(net1),
    .Q(\mod.Arithmetic.CN.I_in[10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _8101_ (.D(\mod.Data_Mem.F_M.out_data[11] ),
    .RN(net2),
    .CLK(net1),
    .Q(\mod.Arithmetic.CN.I_in[11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _8102_ (.D(\mod.Data_Mem.F_M.out_data[12] ),
    .RN(net2),
    .CLK(net1),
    .Q(\mod.Arithmetic.CN.I_in[12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _8103_ (.D(\mod.Data_Mem.F_M.out_data[13] ),
    .RN(net2),
    .CLK(net1),
    .Q(\mod.Arithmetic.CN.I_in[13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _8104_ (.D(\mod.Data_Mem.F_M.out_data[14] ),
    .RN(net2),
    .CLK(net1),
    .Q(\mod.Arithmetic.CN.I_in[14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _8105_ (.D(\mod.Data_Mem.F_M.out_data[15] ),
    .RN(net2),
    .CLK(net1),
    .Q(\mod.Arithmetic.CN.I_in[15] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _8106_ (.D(\mod.Data_Mem.F_M.out_data[16] ),
    .RN(net2),
    .CLK(net1),
    .Q(\mod.Arithmetic.CN.I_in[16] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _8107_ (.D(\mod.Data_Mem.F_M.out_data[17] ),
    .RN(net2),
    .CLK(net1),
    .Q(\mod.Arithmetic.CN.I_in[17] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _8108_ (.D(\mod.Data_Mem.F_M.out_data[18] ),
    .RN(net2),
    .CLK(net1),
    .Q(\mod.Arithmetic.CN.I_in[18] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _8109_ (.D(\mod.Data_Mem.F_M.out_data[19] ),
    .RN(net2),
    .CLK(net1),
    .Q(\mod.Arithmetic.CN.I_in[19] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _8110_ (.D(\mod.Data_Mem.F_M.out_data[20] ),
    .RN(net2),
    .CLK(net1),
    .Q(\mod.Arithmetic.CN.I_in[20] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _8111_ (.D(\mod.Data_Mem.F_M.out_data[21] ),
    .RN(net2),
    .CLK(net1),
    .Q(\mod.Arithmetic.CN.I_in[21] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _8112_ (.D(\mod.Data_Mem.F_M.out_data[22] ),
    .RN(net2),
    .CLK(net1),
    .Q(\mod.Arithmetic.CN.I_in[22] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _8113_ (.D(\mod.Data_Mem.F_M.out_data[23] ),
    .RN(net2),
    .CLK(net1),
    .Q(\mod.Arithmetic.CN.I_in[23] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _8114_ (.D(\mod.Data_Mem.F_M.out_data[24] ),
    .RN(net2),
    .CLK(net1),
    .Q(\mod.Arithmetic.CN.I_in[24] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _8115_ (.D(\mod.Data_Mem.F_M.out_data[25] ),
    .RN(net2),
    .CLK(net1),
    .Q(\mod.Arithmetic.CN.I_in[25] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _8116_ (.D(\mod.Data_Mem.F_M.out_data[26] ),
    .RN(net2),
    .CLK(net1),
    .Q(\mod.Arithmetic.CN.I_in[26] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _8117_ (.D(\mod.Data_Mem.F_M.out_data[27] ),
    .RN(net2),
    .CLK(net1),
    .Q(\mod.Arithmetic.CN.I_in[27] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _8118_ (.D(\mod.Data_Mem.F_M.out_data[28] ),
    .RN(net2),
    .CLK(net1),
    .Q(\mod.Arithmetic.CN.I_in[28] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _8119_ (.D(\mod.Data_Mem.F_M.out_data[29] ),
    .RN(net2),
    .CLK(net1),
    .Q(\mod.Arithmetic.CN.I_in[29] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _8120_ (.D(\mod.Data_Mem.F_M.out_data[30] ),
    .RN(net2),
    .CLK(net1),
    .Q(\mod.Arithmetic.CN.I_in[30] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _8121_ (.D(\mod.Data_Mem.F_M.out_data[31] ),
    .RN(net2),
    .CLK(net1),
    .Q(\mod.Arithmetic.CN.I_in[31] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _8122_ (.D(\mod.Data_Mem.F_M.out_data[32] ),
    .RN(net2),
    .CLK(net1),
    .Q(\mod.Arithmetic.CN.I_in[32] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _8123_ (.D(\mod.Data_Mem.F_M.out_data[33] ),
    .RN(net2),
    .CLK(net1),
    .Q(\mod.Arithmetic.CN.I_in[33] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _8124_ (.D(\mod.Data_Mem.F_M.out_data[34] ),
    .RN(net2),
    .CLK(net1),
    .Q(\mod.Arithmetic.CN.I_in[34] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _8125_ (.D(\mod.Data_Mem.F_M.out_data[35] ),
    .RN(net2),
    .CLK(net1),
    .Q(\mod.Arithmetic.CN.I_in[35] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _8126_ (.D(\mod.Data_Mem.F_M.out_data[36] ),
    .RN(net2),
    .CLK(net1),
    .Q(\mod.Arithmetic.CN.I_in[36] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _8127_ (.D(\mod.Data_Mem.F_M.out_data[37] ),
    .RN(net2),
    .CLK(net1),
    .Q(\mod.Arithmetic.CN.I_in[37] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _8128_ (.D(\mod.Data_Mem.F_M.out_data[38] ),
    .RN(net2),
    .CLK(net1),
    .Q(\mod.Arithmetic.CN.I_in[38] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _8129_ (.D(\mod.Data_Mem.F_M.out_data[39] ),
    .RN(net2),
    .CLK(net1),
    .Q(\mod.Arithmetic.CN.I_in[39] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _8130_ (.D(\mod.Data_Mem.F_M.out_data[40] ),
    .RN(net2),
    .CLK(net1),
    .Q(\mod.Arithmetic.CN.I_in[40] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _8131_ (.D(\mod.Data_Mem.F_M.out_data[41] ),
    .RN(net2),
    .CLK(net1),
    .Q(\mod.Arithmetic.CN.I_in[41] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _8132_ (.D(\mod.Data_Mem.F_M.out_data[42] ),
    .RN(net2),
    .CLK(net1),
    .Q(\mod.Arithmetic.CN.I_in[42] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _8133_ (.D(\mod.Data_Mem.F_M.out_data[43] ),
    .RN(net2),
    .CLK(net1),
    .Q(\mod.Arithmetic.CN.I_in[43] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _8134_ (.D(\mod.Data_Mem.F_M.out_data[44] ),
    .RN(net2),
    .CLK(net1),
    .Q(\mod.Arithmetic.CN.I_in[44] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _8135_ (.D(\mod.Data_Mem.F_M.out_data[45] ),
    .RN(net2),
    .CLK(net1),
    .Q(\mod.Arithmetic.CN.I_in[45] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _8136_ (.D(\mod.Data_Mem.F_M.out_data[46] ),
    .RN(net2),
    .CLK(net1),
    .Q(\mod.Arithmetic.CN.I_in[46] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _8137_ (.D(\mod.Data_Mem.F_M.out_data[47] ),
    .RN(net2),
    .CLK(net1),
    .Q(\mod.Arithmetic.CN.I_in[47] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _8138_ (.D(\mod.Data_Mem.F_M.out_data[48] ),
    .RN(net2),
    .CLK(net1),
    .Q(\mod.Arithmetic.CN.I_in[48] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _8139_ (.D(\mod.Data_Mem.F_M.out_data[49] ),
    .RN(net2),
    .CLK(net1),
    .Q(\mod.Arithmetic.CN.I_in[49] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _8140_ (.D(\mod.Data_Mem.F_M.out_data[50] ),
    .RN(net2),
    .CLK(net1),
    .Q(\mod.Arithmetic.CN.I_in[50] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _8141_ (.D(\mod.Data_Mem.F_M.out_data[51] ),
    .RN(net2),
    .CLK(net1),
    .Q(\mod.Arithmetic.CN.I_in[51] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _8142_ (.D(\mod.Data_Mem.F_M.out_data[52] ),
    .RN(net2),
    .CLK(net1),
    .Q(\mod.Arithmetic.CN.I_in[52] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _8143_ (.D(\mod.Data_Mem.F_M.out_data[53] ),
    .RN(net2),
    .CLK(net1),
    .Q(\mod.Arithmetic.CN.I_in[53] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _8144_ (.D(\mod.Data_Mem.F_M.out_data[54] ),
    .RN(net2),
    .CLK(net1),
    .Q(\mod.Arithmetic.CN.I_in[54] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _8145_ (.D(\mod.Data_Mem.F_M.out_data[55] ),
    .RN(net2),
    .CLK(net1),
    .Q(\mod.Arithmetic.CN.I_in[55] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _8146_ (.D(\mod.Data_Mem.F_M.out_data[56] ),
    .RN(net2),
    .CLK(net1),
    .Q(\mod.Arithmetic.CN.I_in[56] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _8147_ (.D(\mod.Data_Mem.F_M.out_data[57] ),
    .RN(net2),
    .CLK(net1),
    .Q(\mod.Arithmetic.CN.I_in[57] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _8148_ (.D(\mod.Data_Mem.F_M.out_data[58] ),
    .RN(net2),
    .CLK(net1),
    .Q(\mod.Arithmetic.CN.I_in[58] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _8149_ (.D(\mod.Data_Mem.F_M.out_data[59] ),
    .RN(net2),
    .CLK(net1),
    .Q(\mod.Arithmetic.CN.I_in[59] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _8150_ (.D(\mod.Data_Mem.F_M.out_data[60] ),
    .RN(net2),
    .CLK(net1),
    .Q(\mod.Arithmetic.CN.I_in[60] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _8151_ (.D(\mod.Data_Mem.F_M.out_data[61] ),
    .RN(net2),
    .CLK(net1),
    .Q(\mod.Arithmetic.CN.I_in[61] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _8152_ (.D(\mod.Data_Mem.F_M.out_data[62] ),
    .RN(net2),
    .CLK(net1),
    .Q(\mod.Arithmetic.CN.I_in[62] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _8153_ (.D(\mod.Data_Mem.F_M.out_data[63] ),
    .RN(net2),
    .CLK(net1),
    .Q(\mod.Arithmetic.CN.I_in[63] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _8154_ (.D(\mod.Data_Mem.F_M.out_data[64] ),
    .RN(net2),
    .CLK(net1),
    .Q(\mod.Arithmetic.CN.I_in[64] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _8155_ (.D(\mod.Data_Mem.F_M.out_data[65] ),
    .RN(net2),
    .CLK(net1),
    .Q(\mod.Arithmetic.CN.I_in[65] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _8156_ (.D(\mod.Data_Mem.F_M.out_data[66] ),
    .RN(net2),
    .CLK(net1),
    .Q(\mod.Arithmetic.CN.I_in[66] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _8157_ (.D(\mod.Data_Mem.F_M.out_data[67] ),
    .RN(net2),
    .CLK(net1),
    .Q(\mod.Arithmetic.CN.I_in[67] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _8158_ (.D(\mod.Data_Mem.F_M.out_data[68] ),
    .RN(net2),
    .CLK(net1),
    .Q(\mod.Arithmetic.CN.I_in[68] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _8159_ (.D(\mod.Data_Mem.F_M.out_data[69] ),
    .RN(net2),
    .CLK(net1),
    .Q(\mod.Arithmetic.CN.I_in[69] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _8160_ (.D(\mod.Data_Mem.F_M.out_data[70] ),
    .RN(net2),
    .CLK(net1),
    .Q(\mod.Arithmetic.CN.I_in[70] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _8161_ (.D(\mod.Data_Mem.F_M.out_data[71] ),
    .RN(net2),
    .CLK(net1),
    .Q(\mod.Arithmetic.CN.I_in[71] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _8162_ (.D(\mod.Data_Mem.F_M.out_data[72] ),
    .RN(net2),
    .CLK(net1),
    .Q(\mod.Arithmetic.I_out[72] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _8163_ (.D(\mod.Data_Mem.F_M.out_data[73] ),
    .RN(net2),
    .CLK(net1),
    .Q(\mod.Arithmetic.I_out[73] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _8164_ (.D(\mod.Data_Mem.F_M.out_data[74] ),
    .RN(net2),
    .CLK(net1),
    .Q(\mod.Arithmetic.I_out[74] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _8165_ (.D(\mod.Data_Mem.F_M.out_data[75] ),
    .RN(net2),
    .CLK(net1),
    .Q(\mod.Arithmetic.I_out[75] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _8166_ (.D(\mod.Data_Mem.F_M.out_data[76] ),
    .RN(net2),
    .CLK(net1),
    .Q(\mod.Arithmetic.I_out[76] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _8167_ (.D(\mod.Data_Mem.F_M.out_data[77] ),
    .RN(net2),
    .CLK(net1),
    .Q(\mod.Arithmetic.I_out[77] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_2 _8168_ (.D(\mod.Data_Mem.F_M.out_data[78] ),
    .RN(net2),
    .CLK(net1),
    .Q(\mod.Arithmetic.I_out[78] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _8169_ (.D(\mod.Data_Mem.F_M.out_data[79] ),
    .RN(net2),
    .CLK(net1),
    .Q(\mod.Arithmetic.I_out[79] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _8170_ (.D(\mod.P2.dest_reg[0] ),
    .RN(net2),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.dest[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _8171_ (.D(\mod.P2.dest_reg[1] ),
    .RN(net2),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.dest[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _8172_ (.D(\mod.P2.dest_reg[2] ),
    .RN(net2),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.dest[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _8173_ (.D(\mod.P2.dest_reg[4] ),
    .RN(net2),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.dest[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _8174_ (.D(\mod.P2.dest_reg[8] ),
    .RN(net2),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.dest[8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _8175_ (.D(\mod.DM_en ),
    .RN(net2),
    .CLK(net1),
    .Q(\mod.DMen_reg ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _8176_ (.D(\mod.P1.instr_reg[7] ),
    .RN(net2),
    .CLK(net1),
    .Q(\mod.P2.Rout_reg1[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _8177_ (.D(\mod.P1.instr_reg[8] ),
    .RN(net2),
    .CLK(net1),
    .Q(\mod.P2.Rout_reg1[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8178_ (.D(_0288_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.MRAM[3][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8179_ (.D(_0289_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.MRAM[3][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8180_ (.D(_0290_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.MRAM[3][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8181_ (.D(_0291_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.MRAM[3][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8182_ (.D(_0292_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.MRAM[3][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8183_ (.D(_0293_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.MRAM[3][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8184_ (.D(_0294_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.MRAM[3][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8185_ (.D(_0295_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.MRAM[3][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8186_ (.D(_0296_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.MRAM[19][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8187_ (.D(_0297_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.MRAM[19][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8188_ (.D(_0298_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.MRAM[19][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8189_ (.D(_0299_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.MRAM[19][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8190_ (.D(_0300_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.MRAM[19][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8191_ (.D(_0301_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.MRAM[19][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8192_ (.D(_0302_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.MRAM[19][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8193_ (.D(_0303_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.MRAM[19][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _8194_ (.D(net191),
    .RN(net2),
    .CLK(net1),
    .Q(\mod.Arithmetic.CN.F_in[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _8195_ (.D(_0080_),
    .RN(net2),
    .CLK(net1),
    .Q(\mod.I_addr[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _8196_ (.D(_0081_),
    .RN(net2),
    .CLK(net1),
    .Q(\mod.I_addr[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _8197_ (.D(_0082_),
    .RN(net2),
    .CLK(net1),
    .Q(\mod.I_addr[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _8198_ (.D(_0083_),
    .RN(net2),
    .CLK(net1),
    .Q(\mod.I_addr[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _8199_ (.D(_0084_),
    .RN(net2),
    .CLK(net1),
    .Q(\mod.I_addr[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _8200_ (.D(_0085_),
    .RN(net2),
    .CLK(net1),
    .Q(\mod.I_addr[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _8201_ (.D(_0086_),
    .RN(net2),
    .CLK(net1),
    .Q(\mod.I_addr[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _8202_ (.D(_0087_),
    .RN(net2),
    .CLK(net1),
    .Q(\mod.I_addr[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8203_ (.D(_0304_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.MRAM[12][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8204_ (.D(_0305_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.MRAM[12][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8205_ (.D(_0306_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.MRAM[12][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8206_ (.D(_0307_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.MRAM[12][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8207_ (.D(_0308_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.MRAM[12][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8208_ (.D(_0309_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.MRAM[12][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8209_ (.D(_0310_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.MRAM[12][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8210_ (.D(_0311_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.MRAM[12][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8211_ (.D(_0312_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.MRAM[22][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8212_ (.D(_0313_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.MRAM[22][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8213_ (.D(_0314_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.MRAM[22][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8214_ (.D(_0315_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.MRAM[22][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8215_ (.D(_0316_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.MRAM[22][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8216_ (.D(_0317_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.MRAM[22][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8217_ (.D(_0318_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.MRAM[22][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8218_ (.D(_0319_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.MRAM[22][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8219_ (.D(_0320_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.MRAM[29][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8220_ (.D(_0321_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.MRAM[29][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8221_ (.D(_0322_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.MRAM[29][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8222_ (.D(_0323_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.MRAM[29][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8223_ (.D(_0324_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.MRAM[29][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8224_ (.D(_0325_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.MRAM[29][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8225_ (.D(_0326_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.MRAM[29][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8226_ (.D(_0327_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.MRAM[29][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _8227_ (.D(\mod.P1.instr_reg[9] ),
    .RN(net2),
    .CLK(net1),
    .Q(\mod.P2.dest_reg1[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _8228_ (.D(\mod.P1.instr_reg[10] ),
    .RN(net2),
    .CLK(net1),
    .Q(\mod.P2.dest_reg1[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _8229_ (.D(\mod.P1.instr_reg[11] ),
    .RN(net2),
    .CLK(net1),
    .Q(\mod.P2.dest_reg1[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _8230_ (.D(\mod.P1.instr_reg[13] ),
    .RN(net2),
    .CLK(net1),
    .Q(\mod.P2.dest_reg1[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _8231_ (.D(\mod.P1.instr_reg[17] ),
    .RN(net2),
    .CLK(net1),
    .Q(\mod.P2.dest_reg1[8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8232_ (.D(_0328_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.MRAM[2][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8233_ (.D(_0329_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.MRAM[2][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8234_ (.D(_0330_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.MRAM[2][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8235_ (.D(_0331_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.MRAM[2][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8236_ (.D(_0332_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.MRAM[2][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8237_ (.D(_0333_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.MRAM[2][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8238_ (.D(_0334_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.MRAM[2][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8239_ (.D(_0335_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.MRAM[2][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8240_ (.D(_0336_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.MRAM[30][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8241_ (.D(_0337_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.MRAM[30][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8242_ (.D(_0338_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.MRAM[30][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8243_ (.D(_0339_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.MRAM[30][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8244_ (.D(_0340_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.MRAM[30][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8245_ (.D(_0341_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.MRAM[30][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8246_ (.D(_0342_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.MRAM[30][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8247_ (.D(_0343_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.MRAM[30][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8248_ (.D(_0344_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.MRAM[31][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8249_ (.D(_0345_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.MRAM[31][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8250_ (.D(_0346_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.MRAM[31][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8251_ (.D(_0347_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.MRAM[31][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8252_ (.D(_0348_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.MRAM[31][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8253_ (.D(_0349_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.MRAM[31][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8254_ (.D(_0350_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.MRAM[31][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8255_ (.D(_0351_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.MRAM[31][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8256_ (.D(_0352_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.MRAM[5][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8257_ (.D(_0353_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.MRAM[5][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8258_ (.D(_0354_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.MRAM[5][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8259_ (.D(_0355_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.MRAM[5][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8260_ (.D(_0356_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.MRAM[5][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8261_ (.D(_0357_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.MRAM[5][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8262_ (.D(_0358_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.MRAM[5][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8263_ (.D(_0359_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.MRAM[5][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8264_ (.D(_0360_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.MRAM[768][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8265_ (.D(_0361_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.MRAM[768][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8266_ (.D(_0362_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.MRAM[768][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8267_ (.D(_0363_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.MRAM[768][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8268_ (.D(_0364_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.MRAM[768][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8269_ (.D(_0365_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.MRAM[768][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8270_ (.D(_0366_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.MRAM[768][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8271_ (.D(_0367_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.MRAM[768][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8272_ (.D(_0368_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.MRAM[770][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8273_ (.D(_0369_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.MRAM[770][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8274_ (.D(_0370_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.MRAM[770][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8275_ (.D(_0371_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.MRAM[770][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8276_ (.D(_0372_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.MRAM[770][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8277_ (.D(_0373_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.MRAM[770][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8278_ (.D(_0374_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.MRAM[770][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8279_ (.D(_0375_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.MRAM[770][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8280_ (.D(_0376_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.MRAM[771][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8281_ (.D(_0377_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.MRAM[771][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8282_ (.D(_0378_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.MRAM[771][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8283_ (.D(_0379_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.MRAM[771][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8284_ (.D(_0380_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.MRAM[771][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8285_ (.D(_0381_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.MRAM[771][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8286_ (.D(_0382_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.MRAM[771][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8287_ (.D(_0383_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.MRAM[771][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8288_ (.D(_0384_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.MRAM[772][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8289_ (.D(_0385_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.MRAM[772][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8290_ (.D(_0386_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.MRAM[772][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8291_ (.D(_0387_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.MRAM[772][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8292_ (.D(_0388_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.MRAM[772][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8293_ (.D(_0389_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.MRAM[772][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8294_ (.D(_0390_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.MRAM[772][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8295_ (.D(_0391_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.MRAM[772][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8296_ (.D(_0392_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.MRAM[773][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8297_ (.D(_0393_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.MRAM[773][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8298_ (.D(_0394_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.MRAM[773][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8299_ (.D(_0395_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.MRAM[773][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8300_ (.D(_0396_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.MRAM[773][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8301_ (.D(_0397_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.MRAM[773][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8302_ (.D(_0398_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.MRAM[773][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8303_ (.D(_0399_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.MRAM[773][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8304_ (.D(_0400_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.MRAM[774][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8305_ (.D(_0401_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.MRAM[774][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8306_ (.D(_0402_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.MRAM[774][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8307_ (.D(_0403_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.MRAM[774][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8308_ (.D(_0404_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.MRAM[774][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8309_ (.D(_0405_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.MRAM[774][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8310_ (.D(_0406_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.MRAM[774][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8311_ (.D(_0407_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.MRAM[774][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8312_ (.D(_0408_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.MRAM[775][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8313_ (.D(_0409_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.MRAM[775][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8314_ (.D(_0410_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.MRAM[775][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8315_ (.D(_0411_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.MRAM[775][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8316_ (.D(_0412_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.MRAM[775][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8317_ (.D(_0413_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.MRAM[775][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8318_ (.D(_0414_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.MRAM[775][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8319_ (.D(_0415_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.MRAM[775][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8320_ (.D(_0416_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.MRAM[776][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8321_ (.D(_0417_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.MRAM[776][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8322_ (.D(_0418_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.MRAM[776][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8323_ (.D(_0419_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.MRAM[776][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8324_ (.D(_0420_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.MRAM[776][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8325_ (.D(_0421_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.MRAM[776][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8326_ (.D(_0422_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.MRAM[776][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8327_ (.D(_0423_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.MRAM[776][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8328_ (.D(_0424_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.MRAM[777][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8329_ (.D(_0425_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.MRAM[777][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8330_ (.D(_0426_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.MRAM[777][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8331_ (.D(_0427_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.MRAM[777][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8332_ (.D(_0428_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.MRAM[777][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8333_ (.D(_0429_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.MRAM[777][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8334_ (.D(_0430_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.MRAM[777][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8335_ (.D(_0431_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.MRAM[777][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8336_ (.D(_0432_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.MRAM[778][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8337_ (.D(_0433_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.MRAM[778][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8338_ (.D(_0434_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.MRAM[778][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8339_ (.D(_0435_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.MRAM[778][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8340_ (.D(_0436_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.MRAM[778][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8341_ (.D(_0437_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.MRAM[778][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8342_ (.D(_0438_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.MRAM[778][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8343_ (.D(_0439_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.MRAM[778][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8344_ (.D(_0440_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.MRAM[780][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8345_ (.D(_0441_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.MRAM[780][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8346_ (.D(_0442_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.MRAM[780][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8347_ (.D(_0443_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.MRAM[780][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8348_ (.D(_0444_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.MRAM[780][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8349_ (.D(_0445_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.MRAM[780][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8350_ (.D(_0446_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.MRAM[780][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8351_ (.D(_0447_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.MRAM[780][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8352_ (.D(_0448_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.MRAM[781][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8353_ (.D(_0449_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.MRAM[781][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8354_ (.D(_0450_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.MRAM[781][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8355_ (.D(_0451_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.MRAM[781][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8356_ (.D(_0452_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.MRAM[781][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8357_ (.D(_0453_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.MRAM[781][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8358_ (.D(_0454_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.MRAM[781][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8359_ (.D(_0455_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.MRAM[781][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8360_ (.D(_0456_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.MRAM[782][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8361_ (.D(_0457_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.MRAM[782][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8362_ (.D(_0458_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.MRAM[782][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8363_ (.D(_0459_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.MRAM[782][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8364_ (.D(_0460_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.MRAM[782][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8365_ (.D(_0461_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.MRAM[782][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8366_ (.D(_0462_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.MRAM[782][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8367_ (.D(_0463_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.MRAM[782][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8368_ (.D(_0464_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.MRAM[783][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8369_ (.D(_0465_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.MRAM[783][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8370_ (.D(_0466_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.MRAM[783][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8371_ (.D(_0467_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.MRAM[783][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8372_ (.D(_0468_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.MRAM[783][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8373_ (.D(_0469_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.MRAM[783][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8374_ (.D(_0470_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.MRAM[783][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8375_ (.D(_0471_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.MRAM[783][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8376_ (.D(_0472_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.MRAM[784][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8377_ (.D(_0473_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.MRAM[784][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8378_ (.D(_0474_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.MRAM[784][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8379_ (.D(_0475_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.MRAM[784][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8380_ (.D(_0476_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.MRAM[784][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8381_ (.D(_0477_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.MRAM[784][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8382_ (.D(_0478_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.MRAM[784][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8383_ (.D(_0479_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.MRAM[784][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8384_ (.D(_0480_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.MRAM[785][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8385_ (.D(_0481_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.MRAM[785][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8386_ (.D(_0482_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.MRAM[785][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8387_ (.D(_0483_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.MRAM[785][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8388_ (.D(_0484_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.MRAM[785][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8389_ (.D(_0485_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.MRAM[785][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8390_ (.D(_0486_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.MRAM[785][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8391_ (.D(_0487_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.MRAM[785][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8392_ (.D(_0488_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.MRAM[786][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8393_ (.D(_0489_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.MRAM[786][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8394_ (.D(_0490_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.MRAM[786][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8395_ (.D(_0491_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.MRAM[786][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8396_ (.D(_0492_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.MRAM[786][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8397_ (.D(_0493_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.MRAM[786][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8398_ (.D(_0494_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.MRAM[786][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8399_ (.D(_0495_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.MRAM[786][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8400_ (.D(_0496_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.MRAM[787][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8401_ (.D(_0497_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.MRAM[787][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8402_ (.D(_0498_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.MRAM[787][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8403_ (.D(_0499_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.MRAM[787][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8404_ (.D(_0500_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.MRAM[787][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8405_ (.D(_0501_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.MRAM[787][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8406_ (.D(_0502_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.MRAM[787][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8407_ (.D(_0503_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.MRAM[787][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8408_ (.D(_0504_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.MRAM[788][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8409_ (.D(_0505_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.MRAM[788][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8410_ (.D(_0506_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.MRAM[788][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8411_ (.D(_0507_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.MRAM[788][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8412_ (.D(_0508_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.MRAM[788][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8413_ (.D(_0509_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.MRAM[788][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8414_ (.D(_0510_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.MRAM[788][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8415_ (.D(_0511_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.MRAM[788][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8416_ (.D(_0512_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.MRAM[790][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8417_ (.D(_0513_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.MRAM[790][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8418_ (.D(_0514_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.MRAM[790][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8419_ (.D(_0515_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.MRAM[790][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8420_ (.D(_0516_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.MRAM[790][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8421_ (.D(_0517_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.MRAM[790][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8422_ (.D(_0518_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.MRAM[790][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8423_ (.D(_0519_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.MRAM[790][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8424_ (.D(_0520_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.MRAM[791][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8425_ (.D(_0521_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.MRAM[791][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8426_ (.D(_0522_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.MRAM[791][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8427_ (.D(_0523_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.MRAM[791][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8428_ (.D(_0524_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.MRAM[791][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8429_ (.D(_0525_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.MRAM[791][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8430_ (.D(_0526_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.MRAM[791][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8431_ (.D(_0527_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.MRAM[791][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8432_ (.D(_0528_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.MRAM[792][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8433_ (.D(_0529_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.MRAM[792][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8434_ (.D(_0530_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.MRAM[792][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8435_ (.D(_0531_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.MRAM[792][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8436_ (.D(_0532_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.MRAM[792][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8437_ (.D(_0533_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.MRAM[792][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8438_ (.D(_0534_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.MRAM[792][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8439_ (.D(_0535_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.MRAM[792][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8440_ (.D(_0536_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.MRAM[793][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8441_ (.D(_0537_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.MRAM[793][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8442_ (.D(_0538_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.MRAM[793][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8443_ (.D(_0539_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.MRAM[793][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8444_ (.D(_0540_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.MRAM[793][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8445_ (.D(_0541_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.MRAM[793][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8446_ (.D(_0542_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.MRAM[793][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8447_ (.D(_0543_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.MRAM[793][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8448_ (.D(_0544_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.MRAM[794][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8449_ (.D(_0545_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.MRAM[794][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8450_ (.D(_0546_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.MRAM[794][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8451_ (.D(_0547_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.MRAM[794][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8452_ (.D(_0548_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.MRAM[794][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8453_ (.D(_0549_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.MRAM[794][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8454_ (.D(_0550_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.MRAM[794][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8455_ (.D(_0551_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.MRAM[794][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8456_ (.D(_0552_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.MRAM[795][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8457_ (.D(_0553_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.MRAM[795][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8458_ (.D(_0554_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.MRAM[795][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8459_ (.D(_0555_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.MRAM[795][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8460_ (.D(_0556_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.MRAM[795][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8461_ (.D(_0557_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.MRAM[795][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8462_ (.D(_0558_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.MRAM[795][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8463_ (.D(_0559_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.MRAM[795][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8464_ (.D(_0560_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.MRAM[796][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8465_ (.D(_0561_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.MRAM[796][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8466_ (.D(_0562_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.MRAM[796][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8467_ (.D(_0563_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.MRAM[796][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8468_ (.D(_0564_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.MRAM[796][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8469_ (.D(_0565_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.MRAM[796][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8470_ (.D(_0566_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.MRAM[796][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8471_ (.D(_0567_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.MRAM[796][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8472_ (.D(_0568_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.MRAM[797][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8473_ (.D(_0569_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.MRAM[797][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8474_ (.D(_0570_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.MRAM[797][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8475_ (.D(_0571_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.MRAM[797][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8476_ (.D(_0572_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.MRAM[797][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8477_ (.D(_0573_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.MRAM[797][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8478_ (.D(_0574_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.MRAM[797][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8479_ (.D(_0575_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.MRAM[797][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8480_ (.D(_0576_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.MRAM[798][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8481_ (.D(_0577_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.MRAM[798][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8482_ (.D(_0578_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.MRAM[798][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8483_ (.D(_0579_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.MRAM[798][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8484_ (.D(_0580_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.MRAM[798][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8485_ (.D(_0581_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.MRAM[798][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8486_ (.D(_0582_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.MRAM[798][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8487_ (.D(_0583_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.MRAM[798][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8488_ (.D(_0584_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.MRAM[7][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8489_ (.D(_0585_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.MRAM[7][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8490_ (.D(_0586_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.MRAM[7][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8491_ (.D(_0587_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.MRAM[7][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8492_ (.D(_0588_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.MRAM[7][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8493_ (.D(_0589_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.MRAM[7][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8494_ (.D(_0590_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.MRAM[7][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8495_ (.D(_0591_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.MRAM[7][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8496_ (.D(_0000_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.out_data[72] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8497_ (.D(_0001_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.out_data[73] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8498_ (.D(_0002_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.out_data[74] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8499_ (.D(_0003_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.out_data[75] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8500_ (.D(_0004_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.out_data[76] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8501_ (.D(_0005_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.out_data[77] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8502_ (.D(_0006_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.out_data[78] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8503_ (.D(_0007_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.out_data[79] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8504_ (.D(_0008_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.out_data[64] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8505_ (.D(_0009_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.out_data[65] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8506_ (.D(_0010_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.out_data[66] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8507_ (.D(_0011_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.out_data[67] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8508_ (.D(net190),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.out_data[68] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8509_ (.D(net189),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.out_data[69] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8510_ (.D(net188),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.out_data[70] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8511_ (.D(net187),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.out_data[71] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8512_ (.D(_0016_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.out_data[56] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8513_ (.D(_0017_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.out_data[57] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8514_ (.D(_0018_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.out_data[58] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8515_ (.D(_0019_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.out_data[59] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8516_ (.D(net186),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.out_data[60] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8517_ (.D(net185),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.out_data[61] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8518_ (.D(net184),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.out_data[62] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8519_ (.D(net183),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.out_data[63] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8520_ (.D(_0024_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.out_data[48] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8521_ (.D(_0025_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.out_data[49] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8522_ (.D(_0026_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.out_data[50] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8523_ (.D(_0027_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.out_data[51] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8524_ (.D(net182),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.out_data[52] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8525_ (.D(net181),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.out_data[53] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8526_ (.D(net180),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.out_data[54] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8527_ (.D(net179),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.out_data[55] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8528_ (.D(_0032_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.out_data[40] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8529_ (.D(_0033_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.out_data[41] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8530_ (.D(_0034_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.out_data[42] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8531_ (.D(_0035_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.out_data[43] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8532_ (.D(_0036_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.out_data[44] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8533_ (.D(_0037_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.out_data[45] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8534_ (.D(_0038_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.out_data[46] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8535_ (.D(_0039_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.out_data[47] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8536_ (.D(_0040_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.out_data[32] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8537_ (.D(_0041_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.out_data[33] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8538_ (.D(_0042_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.out_data[34] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8539_ (.D(_0043_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.out_data[35] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8540_ (.D(_0044_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.out_data[36] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8541_ (.D(_0045_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.out_data[37] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8542_ (.D(_0046_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.out_data[38] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8543_ (.D(_0047_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.out_data[39] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8544_ (.D(_0048_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.out_data[24] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8545_ (.D(_0049_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.out_data[25] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8546_ (.D(_0050_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.out_data[26] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8547_ (.D(_0051_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.out_data[27] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8548_ (.D(_0052_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.out_data[28] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8549_ (.D(_0053_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.out_data[29] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8550_ (.D(_0054_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.out_data[30] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8551_ (.D(_0055_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.out_data[31] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8552_ (.D(_0056_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.out_data[16] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8553_ (.D(_0057_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.out_data[17] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8554_ (.D(_0058_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.out_data[18] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8555_ (.D(_0059_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.out_data[19] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8556_ (.D(_0060_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.out_data[20] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8557_ (.D(_0061_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.out_data[21] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8558_ (.D(_0062_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.out_data[22] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8559_ (.D(_0063_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.out_data[23] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8560_ (.D(_0064_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.out_data[8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8561_ (.D(_0065_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.out_data[9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8562_ (.D(_0066_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.out_data[10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8563_ (.D(_0067_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.out_data[11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8564_ (.D(_0068_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.out_data[12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8565_ (.D(_0069_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.out_data[13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8566_ (.D(_0070_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.out_data[14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8567_ (.D(_0071_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.out_data[15] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8568_ (.D(_0072_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.out_data[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8569_ (.D(_0073_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.out_data[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8570_ (.D(_0074_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.out_data[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8571_ (.D(_0075_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.out_data[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8572_ (.D(_0076_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.out_data[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8573_ (.D(_0077_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.out_data[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8574_ (.D(_0078_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.out_data[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8575_ (.D(_0079_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.out_data[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8576_ (.D(_0592_),
    .CLK(net1),
    .Q(\mod.Instr_Mem.instruction[8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8577_ (.D(_0593_),
    .CLK(net1),
    .Q(\mod.Instr_Mem.instruction[26] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8578_ (.D(_0594_),
    .CLK(net1),
    .Q(\mod.Instr_Mem.instruction[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8579_ (.D(_0595_),
    .CLK(net1),
    .Q(\mod.Instr_Mem.instruction[13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8580_ (.D(_0596_),
    .CLK(net1),
    .Q(\mod.Instr_Mem.instruction[9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8581_ (.D(_0597_),
    .CLK(net1),
    .Q(\mod.Instr_Mem.instruction[10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8582_ (.D(_0598_),
    .CLK(net1),
    .Q(\mod.Instr_Mem.instruction[22] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8583_ (.D(_0599_),
    .CLK(net1),
    .Q(\mod.Instr_Mem.instruction[23] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8584_ (.D(_0600_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.MRAM[9][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8585_ (.D(_0601_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.MRAM[9][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8586_ (.D(_0602_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.MRAM[9][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8587_ (.D(_0603_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.MRAM[9][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8588_ (.D(_0604_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.MRAM[9][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8589_ (.D(_0605_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.MRAM[9][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8590_ (.D(_0606_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.MRAM[9][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8591_ (.D(_0607_),
    .CLK(net1),
    .Q(\mod.Data_Mem.F_M.MRAM[9][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8592_ (.D(_0608_),
    .CLK(net1),
    .Q(\mod.Instr_Mem.instruction[11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8593_ (.D(_0609_),
    .CLK(net1),
    .Q(\mod.Instr_Mem.instruction[17] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8594_ (.D(_0610_),
    .CLK(net1),
    .Q(\mod.Instr_Mem.instruction[24] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8595_ (.D(_0611_),
    .CLK(net1),
    .Q(\mod.Instr_Mem.instruction[30] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8498__D (.I(_0002_));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_12 (.ZN(net12));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_13 (.ZN(net13));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_14 (.ZN(net14));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_15 (.ZN(net15));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_16 (.ZN(net16));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_17 (.ZN(net17));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_18 (.ZN(net18));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_19 (.ZN(net19));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_20 (.ZN(net20));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_21 (.ZN(net21));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_22 (.ZN(net22));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_23 (.ZN(net23));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_24 (.ZN(net24));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_25 (.ZN(net25));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_26 (.ZN(net26));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_27 (.ZN(net27));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_28 (.ZN(net28));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_29 (.ZN(net29));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_30 (.ZN(net30));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_31 (.ZN(net31));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_32 (.ZN(net32));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_33 (.ZN(net33));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_34 (.ZN(net34));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_35 (.ZN(net35));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_36 (.ZN(net36));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_37 (.ZN(net37));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_38 (.ZN(net38));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_39 (.ZN(net39));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_40 (.ZN(net40));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_41 (.ZN(net41));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_42 (.ZN(net42));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_43 (.ZN(net43));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_44 (.ZN(net44));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_45 (.ZN(net45));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_46 (.ZN(net46));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_47 (.ZN(net47));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_48 (.ZN(net48));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_49 (.ZN(net49));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_50 (.ZN(net50));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_51 (.ZN(net51));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_52 (.ZN(net52));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_53 (.ZN(net53));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_54 (.ZN(net54));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_55 (.ZN(net55));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_56 (.ZN(net56));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_57 (.ZN(net57));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_58 (.ZN(net58));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_59 (.ZN(net59));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_60 (.ZN(net60));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_61 (.ZN(net61));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_62 (.ZN(net62));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_63 (.ZN(net63));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_64 (.ZN(net64));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_65 (.ZN(net65));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_66 (.ZN(net66));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_67 (.ZN(net67));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_68 (.ZN(net68));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_69 (.ZN(net69));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_70 (.ZN(net70));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_71 (.ZN(net71));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_72 (.ZN(net72));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_73 (.ZN(net73));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_74 (.ZN(net74));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_75 (.ZN(net75));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_76 (.ZN(net76));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_77 (.ZN(net77));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_78 (.ZN(net78));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_79 (.ZN(net79));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_80 (.ZN(net80));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_81 (.ZN(net81));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_82 (.ZN(net82));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_83 (.ZN(net83));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_84 (.ZN(net84));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_85 (.ZN(net85));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_86 (.ZN(net86));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_87 (.ZN(net87));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_88 (.ZN(net88));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_89 (.ZN(net89));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_90 (.ZN(net90));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_91 (.ZN(net91));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_92 (.ZN(net92));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_93 (.ZN(net93));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_94 (.ZN(net94));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_95 (.ZN(net95));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_96 (.ZN(net96));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_97 (.ZN(net97));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_98 (.ZN(net98));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_99 (.ZN(net99));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_100 (.ZN(net100));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_101 (.ZN(net101));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_102 (.ZN(net102));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_103 (.ZN(net103));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_104 (.ZN(net104));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_105 (.ZN(net105));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_106 (.ZN(net106));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_107 (.ZN(net107));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_108 (.ZN(net108));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_109 (.ZN(net109));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_110 (.ZN(net110));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_111 (.ZN(net111));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_112 (.ZN(net112));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_113 (.ZN(net113));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_114 (.ZN(net114));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_115 (.ZN(net115));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_116 (.ZN(net116));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_117 (.ZN(net117));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_118 (.ZN(net118));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_119 (.ZN(net119));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_120 (.ZN(net120));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_121 (.ZN(net121));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_122 (.ZN(net122));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_123 (.ZN(net123));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_124 (.ZN(net124));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_125 (.ZN(net125));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_126 (.ZN(net126));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_127 (.ZN(net127));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_128 (.ZN(net128));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_129 (.ZN(net129));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_130 (.ZN(net130));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_131 (.ZN(net131));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_132 (.ZN(net132));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_133 (.ZN(net133));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_134 (.ZN(net134));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_135 (.ZN(net135));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_136 (.ZN(net136));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_137 (.ZN(net137));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_138 (.ZN(net138));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_139 (.ZN(net139));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_140 (.ZN(net140));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_141 (.ZN(net141));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_142 (.ZN(net142));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_143 (.ZN(net143));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_144 (.ZN(net144));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_145 (.ZN(net145));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_146 (.ZN(net146));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_147 (.ZN(net147));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_148 (.ZN(net148));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_149 (.ZN(net149));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_150 (.ZN(net150));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_151 (.ZN(net151));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_152 (.ZN(net152));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_153 (.ZN(net153));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_154 (.ZN(net154));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_155 (.ZN(net155));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_156 (.ZN(net156));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_157 (.ZN(net157));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_158 (.ZN(net158));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_159 (.ZN(net159));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_160 (.ZN(net160));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_161 (.ZN(net161));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_162 (.ZN(net162));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_163 (.ZN(net163));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_164 (.ZN(net164));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_165 (.ZN(net165));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_166 (.ZN(net166));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_167 (.ZN(net167));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_168 (.ZN(net168));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_169 (.ZN(net169));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_170 (.ZN(net170));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_171 (.ZN(net171));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_172 (.ZN(net172));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_173 (.ZN(net173));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_174 (.ZN(net174));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_175 (.ZN(net175));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_176 (.ZN(net176));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_177 (.ZN(net177));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_178 (.ZN(net178));
 gf180mcu_fd_sc_mcu7t5v0__tiel _8527__179 (.ZN(net179));
 gf180mcu_fd_sc_mcu7t5v0__tiel _8526__180 (.ZN(net180));
 gf180mcu_fd_sc_mcu7t5v0__tiel _8525__181 (.ZN(net181));
 gf180mcu_fd_sc_mcu7t5v0__tiel _8524__182 (.ZN(net182));
 gf180mcu_fd_sc_mcu7t5v0__tiel _8519__183 (.ZN(net183));
 gf180mcu_fd_sc_mcu7t5v0__tiel _8518__184 (.ZN(net184));
 gf180mcu_fd_sc_mcu7t5v0__tiel _8517__185 (.ZN(net185));
 gf180mcu_fd_sc_mcu7t5v0__tiel _8516__186 (.ZN(net186));
 gf180mcu_fd_sc_mcu7t5v0__tiel _8511__187 (.ZN(net187));
 gf180mcu_fd_sc_mcu7t5v0__tiel _8510__188 (.ZN(net188));
 gf180mcu_fd_sc_mcu7t5v0__tiel _8509__189 (.ZN(net189));
 gf180mcu_fd_sc_mcu7t5v0__tiel _8508__190 (.ZN(net190));
 gf180mcu_fd_sc_mcu7t5v0__tieh _8194__191 (.Z(net191));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_0 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_6 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_7 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_8 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_9 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_10 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_11 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_12 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_13 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_14 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_15 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_16 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_17 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_18 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_19 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_20 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_21 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_22 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_23 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_24 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_25 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_26 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_27 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_28 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_29 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_30 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_31 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_32 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_33 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_34 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_35 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_36 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_37 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_38 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_39 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_40 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_41 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_42 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_43 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_44 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_45 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_46 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_47 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_48 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_49 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_50 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_51 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_52 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_53 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_54 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_55 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_56 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_57 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_58 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_59 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_60 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_61 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_62 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_63 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_64 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_65 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_66 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_67 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_68 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_69 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_70 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_71 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_72 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_73 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_74 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_75 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_76 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_77 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_78 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_79 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_80 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_81 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_82 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_83 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_84 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_85 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_86 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_87 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_88 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_89 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_90 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_91 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_92 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_93 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_94 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_95 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_96 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_97 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_98 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_99 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_100 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_101 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_102 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_103 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_104 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_105 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_106 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_107 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_108 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_109 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_110 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_111 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_112 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_113 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_114 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_115 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_116 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_117 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_118 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_119 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_120 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_121 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_122 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_123 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_124 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_125 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_126 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_127 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_128 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_129 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_130 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_131 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_132 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_133 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_134 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_135 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_136 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_137 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_138 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_139 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_140 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_141 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_142 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_143 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_144 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_145 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_146 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_147 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_148 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_149 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_150 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_151 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_152 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_153 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_154 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_155 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_156 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_157 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_158 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_159 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_160 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_161 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_162 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_163 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_164 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_165 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_166 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_167 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_168 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_169 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_170 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_171 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_172 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_173 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_174 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_175 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_176 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_177 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_178 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_179 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_180 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_181 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_182 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_183 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_184 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_185 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_186 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_187 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_188 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_189 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_190 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_191 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_192 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_193 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_194 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_195 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_196 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_197 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_198 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_199 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_200 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_201 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_202 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_203 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_204 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_205 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_206 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_207 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_208 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_209 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_210 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_211 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_212 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_213 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_214 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_215 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_216 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_217 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_218 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_219 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_220 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_221 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_222 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_223 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_224 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_225 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_226 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_227 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_228 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_229 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_230 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_231 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_232 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_233 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_234 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_235 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_236 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_237 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_238 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_239 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_240 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_241 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_242 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_243 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_244 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_245 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_246 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_247 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_248 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_249 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_250 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_251 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_252 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_253 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_254 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_255 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_256 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_257 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_258 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_259 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_260 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_261 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_262 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_263 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_264 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_265 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_266 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_267 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_268 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_269 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_270 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_271 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_272 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_273 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_274 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_275 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_276 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_277 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_278 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_279 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_280 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_281 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_282 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_283 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_284 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_285 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_286 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_287 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_288 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_289 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_290 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_291 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_292 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_293 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_294 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_295 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_296 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_297 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_298 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_299 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_300 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_301 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_302 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_303 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_304 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_305 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_306 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_307 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_308 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_309 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_310 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_311 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_312 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_313 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_314 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_315 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_316 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_317 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_318 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_319 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_320 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_321 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_322 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_323 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_324 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_325 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_326 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_327 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_328 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_329 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_330 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_331 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_332 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_333 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_334 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_335 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_336 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_337 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_338 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_339 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_340 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_341 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_342 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_343 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_344 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_345 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_346 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_347 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_348 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_349 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_350 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_351 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_352 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_353 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_354 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_355 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_356 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_357 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_358 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_359 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_360 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_361 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_362 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_363 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_364 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_365 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_366 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_367 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_368 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_369 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_370 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_371 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_372 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_373 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_374 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_375 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_376 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_377 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_378 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_379 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_380 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_381 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_382 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_383 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_384 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_385 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_386 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_387 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_388 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_389 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_390 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_391 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_392 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_393 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_394 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_395 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_396 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_397 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_398 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_399 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_400 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_401 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_402 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_403 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_404 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_405 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_406 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_407 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_408 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_409 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_410 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_411 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_412 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_413 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_414 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_415 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_416 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_417 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_418 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_419 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_420 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_421 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_422 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_423 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_424 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_425 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_426 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_427 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_428 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_429 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_430 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_431 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_432 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_433 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_434 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_435 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_436 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_437 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_438 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_439 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_440 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_441 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_442 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_443 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_444 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_445 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_446 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_447 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_448 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_449 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_450 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_451 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_452 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_453 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_454 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_455 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_456 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_457 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_458 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_459 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_460 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_461 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_462 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_463 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_464 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_465 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_466 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_467 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_468 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_469 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_470 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_471 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_472 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_473 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_474 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_475 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_476 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_477 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_478 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_479 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_480 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_481 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_482 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_483 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_484 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_485 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_486 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_487 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_488 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_489 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_490 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_491 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_492 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_493 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_494 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_495 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_496 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_497 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_498 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_499 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_500 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_501 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_502 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_503 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_504 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_505 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_506 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_507 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_508 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_509 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_510 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_511 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_512 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_513 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_514 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_515 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_516 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_517 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_518 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_519 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_520 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_521 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_522 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_523 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_524 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_525 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_526 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_527 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_528 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_529 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_530 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_531 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_532 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_533 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_534 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_535 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_536 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_537 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_538 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_539 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_540 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_541 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_542 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_543 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_544 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_545 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_546 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_547 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_548 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_549 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_550 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_551 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_552 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_553 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_554 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_555 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_556 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_557 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_558 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_559 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_560 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_561 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_562 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_563 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_564 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_565 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_566 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_567 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_568 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_569 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_570 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_571 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_572 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_573 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_574 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_575 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_576 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_577 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_578 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_579 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_580 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_581 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_582 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_583 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_584 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_585 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_586 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_587 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_588 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_589 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_590 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_591 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_592 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_593 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_594 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_595 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_596 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_597 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_598 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_599 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_600 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_601 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_602 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_603 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_604 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_605 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_606 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_607 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_608 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_609 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_610 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_611 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_612 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_613 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_614 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_615 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_616 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_617 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_618 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_619 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_620 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_621 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_622 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_623 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_624 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_625 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_626 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_627 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_628 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_629 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_630 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_631 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_632 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_633 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_634 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_635 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_636 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_637 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_638 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_639 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_640 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_641 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_642 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_643 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_644 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_645 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_646 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_647 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_648 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_649 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_650 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_651 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_652 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_653 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_654 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_655 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_656 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_657 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_658 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_659 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_660 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_661 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_662 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_663 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_664 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_665 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_666 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_667 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_668 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_669 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_670 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_671 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_672 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_673 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_674 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_675 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_676 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_677 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_678 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_679 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_680 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_681 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_682 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_683 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_684 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_685 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_686 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_687 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_688 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_689 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_690 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_691 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_692 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_693 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_694 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_695 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_696 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_697 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_698 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_699 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_700 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_701 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_702 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_703 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_704 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_705 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_706 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_707 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_708 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_709 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_710 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_711 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_712 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_713 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_714 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_715 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_716 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_717 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_718 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_719 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_720 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_721 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_722 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_723 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_724 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_725 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_726 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_727 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_728 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_729 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_730 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_731 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_732 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_733 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_734 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_735 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_736 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_737 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_738 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_739 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_740 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_741 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_742 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_743 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_744 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_745 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_746 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_747 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_748 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_749 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_750 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_751 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_752 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_753 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_754 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_755 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_756 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_757 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_758 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_759 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_760 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_761 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_762 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_763 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_764 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_765 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_766 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_767 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_768 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_769 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_770 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_771 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_772 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_773 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_774 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_775 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_776 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_777 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_778 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_779 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_780 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_781 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_782 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_783 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_784 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_785 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_786 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_787 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_788 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_789 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_790 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_791 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_792 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_793 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_794 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_795 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_796 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_797 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_798 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_799 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_800 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_801 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_802 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_803 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_804 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_805 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_806 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_807 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_808 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_809 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_810 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_811 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_812 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_813 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_814 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_815 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_816 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_817 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_818 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_819 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_820 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_821 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_822 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_823 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_824 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_825 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_826 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_827 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_828 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_829 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_830 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_831 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_832 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_833 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_834 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_835 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_836 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_837 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_838 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_839 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_840 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_841 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_842 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_843 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_844 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_845 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_846 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_847 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_848 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_849 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_850 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_851 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_852 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_853 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_854 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_855 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_856 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_857 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_858 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_859 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_860 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_861 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_862 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_863 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_864 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_865 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_866 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_867 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_868 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_869 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_870 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_871 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_872 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_873 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_874 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_875 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_876 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_877 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_878 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_879 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_880 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_881 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_882 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_883 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_884 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_885 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_886 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_887 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_888 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_889 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_890 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_891 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_892 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_893 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_894 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_895 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_896 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_897 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_898 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_899 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_900 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_901 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_902 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_903 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_904 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_905 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_906 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_907 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_908 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_909 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_910 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_911 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_912 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_913 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_914 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_915 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_916 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_917 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_918 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_919 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_920 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_921 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_922 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_923 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_924 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_925 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_926 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_927 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_928 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_929 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_930 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_931 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_932 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_933 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_934 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_935 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_936 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_937 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_938 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_939 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_940 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_941 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_942 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_943 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_944 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_945 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_946 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_947 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_948 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_949 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_950 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_951 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_952 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_953 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_954 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_955 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_956 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_957 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_958 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_959 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_960 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_961 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_962 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_963 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_964 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_965 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_966 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_967 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_968 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_969 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_970 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_971 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_972 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_973 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_974 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_975 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_976 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_977 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_978 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_979 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_980 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_981 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_982 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_983 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_984 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_985 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_986 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_987 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_988 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_989 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_990 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_991 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_992 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_993 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_994 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_995 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_996 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_997 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_998 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_999 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1000 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1016 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1018 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1020 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1029 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1030 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1032 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1035 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1050 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1051 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1053 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1055 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1057 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1058 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1059 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1065 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1066 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1068 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1069 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1071 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1072 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1073 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1075 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1077 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1080 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1085 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1088 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1089 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1090 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1092 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1093 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1094 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1100 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1101 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1103 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1104 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1107 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1108 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1110 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1114 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1120 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1121 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1123 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1124 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1125 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1127 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1128 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1129 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1136 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1137 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1139 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1140 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1142 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1143 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1144 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1146 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1148 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1155 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1156 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1158 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1159 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1160 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1162 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1163 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1164 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1167 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1171 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1172 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1175 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1178 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1179 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1181 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1182 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1185 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1187 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1190 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1191 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1193 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1194 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1195 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1196 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1197 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1198 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1199 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1201 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1203 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1207 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1208 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1210 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1211 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1213 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1214 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1215 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1219 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1225 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1226 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1228 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1229 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1230 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1231 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1232 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1233 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1234 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1235 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1236 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1238 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1240 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1242 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1243 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1245 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1246 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1247 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1248 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1249 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1250 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1252 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1253 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1254 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1255 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1258 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1260 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1261 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1263 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1264 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1265 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1266 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1267 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1268 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1269 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1270 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1271 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1272 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1274 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1275 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1278 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1279 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1281 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1282 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1283 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1284 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1285 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1286 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1287 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1288 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1289 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1290 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1292 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1293 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1295 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1296 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1298 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1299 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1300 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1301 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1302 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1303 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1304 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1305 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1306 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1307 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1309 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1310 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1311 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1313 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1314 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1316 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1317 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1318 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1319 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1320 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1321 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1322 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1323 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1324 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1325 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1327 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1328 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1329 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1330 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1331 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1333 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1334 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1335 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1336 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1337 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1338 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1339 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1340 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1341 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1342 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1343 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1345 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1346 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1349 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1350 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1352 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1353 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1354 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1355 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1356 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1357 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1358 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1359 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1360 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1362 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1364 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1365 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1366 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1368 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1369 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1370 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1371 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1372 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1373 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1374 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1375 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1376 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1377 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1378 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1380 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1381 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1382 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1384 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1385 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1387 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1388 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1389 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1390 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1391 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1392 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1393 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1394 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1395 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1397 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1398 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1400 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1401 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1403 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1404 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1405 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1406 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1407 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1408 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1409 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1410 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1411 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1412 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1413 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1414 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1416 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1417 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1418 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1420 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1421 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1423 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1424 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1425 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1426 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1427 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1428 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1429 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1430 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1432 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1433 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1434 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1435 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1436 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1438 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1439 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1440 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1441 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1442 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1443 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1444 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1445 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1446 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1447 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1448 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1449 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1451 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1452 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1453 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1455 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1456 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1458 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1459 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1460 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1461 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1462 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1463 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1464 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1465 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1467 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1468 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1469 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1470 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1471 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1473 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1474 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1475 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1476 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1477 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1478 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1479 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1480 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1481 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1482 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1483 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1484 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1485 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1487 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1488 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1489 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1491 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1492 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1494 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1495 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1496 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1497 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1498 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1499 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1500 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1502 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1503 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1504 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1505 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1506 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1508 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1509 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1510 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1511 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1512 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1513 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1514 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1515 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1516 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1517 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1518 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1519 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1520 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1522 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1523 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1524 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1526 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1527 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1529 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1530 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1531 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1532 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1533 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1534 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1535 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1537 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1538 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1539 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1540 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1541 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1543 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1544 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1545 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1546 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1547 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1548 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1549 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1550 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1551 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1552 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1553 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1554 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1555 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1556 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1558 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1559 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1562 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1563 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1565 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1566 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1567 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1568 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1569 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1570 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1572 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1573 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1574 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1575 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1578 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1579 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1581 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1582 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1583 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1584 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1585 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1586 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1587 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1588 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1589 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1590 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1591 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1593 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1594 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1595 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1597 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1598 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1600 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1601 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1602 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1603 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1604 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1605 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1607 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1608 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1609 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1610 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1611 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1613 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1614 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1615 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1616 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1617 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1618 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1619 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1620 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1621 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1622 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1623 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1624 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1625 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1626 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1627 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1629 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1630 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1631 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1633 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1634 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1636 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1637 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1638 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1639 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1640 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1642 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1643 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1644 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1645 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1646 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1648 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1649 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1650 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1651 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1652 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1653 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1654 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1655 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1656 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1657 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1658 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1659 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1660 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1661 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1662 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1664 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1665 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1666 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1668 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1669 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1671 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1672 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1673 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1674 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1675 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1677 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1678 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1679 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1680 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1681 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1683 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1684 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1685 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1686 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1687 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1688 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1689 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1690 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1691 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1692 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1693 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1694 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1695 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1696 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1697 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1698 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1700 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1701 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1702 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1704 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1705 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1707 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1708 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1709 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1710 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1712 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1713 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1714 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1715 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1716 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1718 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1719 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1720 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1721 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1722 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1723 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1724 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1725 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1726 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1727 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1728 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1729 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1730 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1731 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1732 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1733 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1735 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1736 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1737 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1739 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1740 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1742 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1743 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1744 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1745 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1747 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1748 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1749 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1750 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1751 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1753 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1755 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1756 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1759 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1760 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1761 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1762 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1763 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1764 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1765 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1766 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1767 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1768 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1769 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1771 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1772 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1773 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1775 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1776 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1778 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1779 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1780 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1781 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1782 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1783 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1784 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1785 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1786 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1787 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1788 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1789 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1790 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1791 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1792 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1793 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1794 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1795 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1796 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1797 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1798 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1799 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1800 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1801 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1802 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1803 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1804 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1806 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1807 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1808 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1810 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1811 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1813 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1814 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1815 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1816 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1817 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1818 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1819 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1820 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1821 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1822 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1823 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1824 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1825 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1826 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1827 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1828 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1829 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1830 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1831 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1832 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1833 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1834 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1835 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1836 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1837 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1838 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1839 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1840 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1842 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1843 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1844 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1846 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1847 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1849 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1850 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1851 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1852 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1853 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1854 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1855 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1856 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1857 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1858 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1859 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1860 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1861 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1862 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1863 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1864 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1865 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1866 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1867 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1868 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1869 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1870 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1871 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1872 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1873 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1874 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1875 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1877 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1878 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1879 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1881 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1882 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1884 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1885 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1886 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1887 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1888 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1889 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1890 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1891 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1892 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1893 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1894 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1895 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1896 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1897 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1898 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1899 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1900 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1901 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1902 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1903 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1904 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1905 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1906 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1907 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1908 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1909 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1910 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1911 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1913 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1914 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1915 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1917 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1918 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1920 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1921 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1922 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1923 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1924 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1925 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1926 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1927 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1928 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1929 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1930 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1931 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1932 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1933 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1934 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1936 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1938 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1939 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1940 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1941 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1942 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1943 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1944 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1945 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1946 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1947 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1948 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1949 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1950 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1951 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1952 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1953 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1954 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1955 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1956 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1957 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1958 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1959 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1960 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1961 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1962 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1963 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1964 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1965 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1966 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1967 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1968 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1969 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1970 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1971 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1972 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1973 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1974 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1975 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1976 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1977 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1978 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1979 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1980 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1981 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1982 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1983 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1984 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1985 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1986 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1987 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1988 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1989 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1990 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1991 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1992 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1993 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1994 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1995 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1996 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1997 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1998 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1999 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2000 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2001 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2002 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2003 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2004 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2005 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2006 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2007 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2008 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2009 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2010 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2011 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2012 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2013 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2014 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2015 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2016 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2017 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2018 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2019 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2020 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2021 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2022 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2023 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2024 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2025 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2026 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2027 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2028 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2029 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2030 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2031 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2032 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2033 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2034 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2035 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2036 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2037 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2038 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2039 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2040 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2041 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2042 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2043 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2044 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2045 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2046 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2047 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2048 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2049 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2050 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2051 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2052 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2053 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2054 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2055 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2056 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2057 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2058 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2059 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2060 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2061 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2062 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2063 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2064 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2065 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2066 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2067 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2068 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2069 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2070 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2071 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2072 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2073 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2074 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2075 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2076 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2077 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2078 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2079 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2080 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2081 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2082 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2083 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2084 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2085 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2086 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2087 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2088 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2089 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2090 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2091 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2092 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2093 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2094 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2095 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2096 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2097 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2098 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2099 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2100 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2101 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2102 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2103 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2104 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2105 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2106 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2107 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2108 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2109 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2110 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2111 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2112 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2113 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2114 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2115 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2116 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2117 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2118 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2119 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2120 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2121 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2122 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2123 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2124 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2125 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2126 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2127 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2128 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2129 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2130 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2132 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2133 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2134 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2135 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2136 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2137 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2138 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2139 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2140 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2141 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2142 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2143 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2144 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2145 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2146 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2147 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2148 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2149 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2150 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2151 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2152 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2153 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2154 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2155 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2156 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2157 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2158 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2159 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2160 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2161 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2162 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2163 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2164 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2165 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2166 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2167 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2168 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2169 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2170 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2171 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2172 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2173 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2174 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2175 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2176 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2177 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2178 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2179 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2180 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2181 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2182 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2183 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2184 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2185 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2186 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2187 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2188 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2189 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2190 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2191 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2192 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2193 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2194 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2195 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2196 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2197 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2198 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2199 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2200 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2201 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2202 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2203 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2204 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2205 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2206 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2207 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2208 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2209 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2210 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2211 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2212 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2213 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2214 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2215 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2216 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2217 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2218 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2219 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2220 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2221 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2222 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2223 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2224 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2225 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2226 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2227 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2228 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2229 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2230 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2231 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2232 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2233 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2234 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2235 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2236 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2237 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2238 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2239 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2240 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2241 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2242 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2243 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2244 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2245 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2246 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2247 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2248 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2249 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2250 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2251 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2252 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2253 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2254 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2255 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2256 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2257 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2258 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2259 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2260 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2261 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2262 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2263 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2264 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2265 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2266 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2267 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2268 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2269 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2270 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2271 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2272 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2273 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2274 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2275 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2276 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2277 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2278 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2279 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2280 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2281 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2282 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2283 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2284 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2285 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2286 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2287 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2288 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2289 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2290 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2291 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2292 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2293 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2294 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2295 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2296 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2297 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2298 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2299 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2300 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2301 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2302 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2303 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2304 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2305 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2306 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2307 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2308 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2309 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2310 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2311 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2312 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2313 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2314 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2315 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2316 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2317 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2318 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2319 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2320 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2321 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2322 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2323 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2324 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2325 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2326 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2327 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2328 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2329 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2330 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2331 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2332 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2333 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2334 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2335 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2336 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2337 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2338 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2339 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2340 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2341 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2342 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2343 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2344 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2345 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2346 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2347 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2348 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2349 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2350 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2351 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2352 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2353 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2354 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2355 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2356 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2357 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2358 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2359 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2360 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2361 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2362 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2363 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2364 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2365 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2366 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2367 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2368 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2369 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2370 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2371 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2372 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2373 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2374 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2375 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2376 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2377 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2378 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2379 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2380 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2381 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2382 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2383 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2384 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2385 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2386 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2387 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2388 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2389 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2390 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2391 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2392 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2393 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2394 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2395 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2396 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2397 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2398 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2399 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2400 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2401 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2402 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2403 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2404 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2405 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2406 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2407 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2408 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2409 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2410 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2411 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2412 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2413 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2414 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2415 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2416 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2417 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2418 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2419 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2420 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2421 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2422 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2423 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2424 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2425 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2426 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2427 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2428 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2429 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2430 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2431 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2432 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2433 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2434 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2435 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2436 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2437 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2438 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2439 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2440 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2441 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2442 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2443 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2444 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2445 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2446 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2447 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2448 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2449 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2450 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2451 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2452 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2453 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2454 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2455 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2456 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2457 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2458 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2459 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2460 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2461 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2462 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2463 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2464 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2465 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2466 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2467 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2468 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2469 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2470 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2471 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2472 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2473 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2474 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2475 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2476 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2477 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2478 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2479 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2480 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2481 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2482 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2483 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2484 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2485 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2486 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2487 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2488 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2489 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2490 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2491 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2492 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2493 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2494 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2495 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2496 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2497 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2498 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2499 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2500 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2501 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2502 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2503 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2504 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2505 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2506 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2507 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2508 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2509 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2510 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2511 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2512 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2513 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2514 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2515 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2516 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2517 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2518 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2519 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2520 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2521 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2522 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2523 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2524 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2525 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2526 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2527 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2528 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2529 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2530 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2531 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2532 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2533 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2534 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2535 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2536 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2537 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2538 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2539 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2540 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2541 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2542 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2543 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2544 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2545 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2546 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2547 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2548 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2549 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2550 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2551 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2552 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2553 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2554 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2555 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2556 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2557 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2558 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2559 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2560 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2561 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2562 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2563 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2564 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2565 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2566 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2567 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2568 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2569 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2570 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2571 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2572 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2573 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2574 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2575 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2576 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2577 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2578 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2579 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2580 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2581 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2582 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2583 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2584 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2585 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2586 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2587 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2588 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2589 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2590 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2591 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2592 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2593 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2594 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2595 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2596 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2597 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2598 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2599 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2600 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2601 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2602 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2603 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2604 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2605 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2606 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2607 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2608 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2609 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2610 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2611 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2612 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2613 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2614 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2615 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2616 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2617 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2618 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2619 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2620 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2621 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2622 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2623 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2624 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2625 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2626 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2627 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2628 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2629 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2630 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2631 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2632 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2633 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2634 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2635 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2636 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2637 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2638 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2639 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2640 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2641 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2642 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2643 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2644 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2645 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2646 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2647 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2648 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2649 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2650 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2651 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2652 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2653 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2654 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2655 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2656 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2657 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2658 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2659 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2660 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2661 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2662 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2663 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2664 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2665 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2666 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2667 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2668 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2669 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2670 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2671 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2672 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2673 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2674 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2675 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2676 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2677 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2678 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2679 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2680 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2681 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2682 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2683 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2684 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2685 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2686 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2687 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2688 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2689 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2690 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2691 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2692 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2693 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2694 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2695 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2696 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2697 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2698 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2699 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2700 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2701 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2702 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2703 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2704 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2705 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2706 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2707 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2708 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2709 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2710 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2711 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2712 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2713 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2714 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2715 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2716 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2717 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2718 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2719 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2720 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2721 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2722 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2723 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2724 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2725 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2726 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2727 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2728 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2729 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2730 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2731 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2732 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2733 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2734 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2735 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2736 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2737 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2738 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2739 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2740 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2741 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2742 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2743 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2744 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2745 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2746 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2747 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2748 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2749 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2750 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2751 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2752 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2753 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2754 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2755 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2756 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2757 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2758 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2759 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2760 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2761 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2762 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2763 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2764 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2765 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2766 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2767 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2768 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2769 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2770 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2771 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2772 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2773 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2774 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2775 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2776 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2777 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2778 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2779 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2780 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2781 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2782 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2783 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2784 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2785 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2786 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2787 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2788 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2789 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2790 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2791 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2792 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2793 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2794 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2795 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2796 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2797 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2798 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2799 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2800 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2801 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2802 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2803 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2804 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2805 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2806 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2807 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2808 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2809 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2810 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2811 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2812 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2813 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2814 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2815 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2816 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2817 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2818 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2819 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2820 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2821 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2822 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2823 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2824 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2825 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2826 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2827 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2828 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2829 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2830 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2831 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2832 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2833 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2834 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2835 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2836 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2837 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2838 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2839 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2840 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2841 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2842 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2843 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2844 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2845 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2846 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2847 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2848 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2849 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2850 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2851 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2852 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2853 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2854 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2855 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2856 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2857 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2858 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2859 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2860 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2861 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2862 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2863 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2864 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2865 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2866 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2867 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2868 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2869 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2870 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2871 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2872 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2873 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2874 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2875 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2876 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2877 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2878 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2879 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2880 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2881 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2882 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2883 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2884 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2885 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2886 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2887 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2888 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2889 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2890 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2891 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2892 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2893 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2894 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2895 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2896 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2897 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2898 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2899 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2900 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2901 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2902 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2903 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2904 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2905 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2906 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2907 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2908 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2909 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2910 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2911 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2912 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2913 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2914 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2915 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2916 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2917 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2918 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2919 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2920 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2921 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2922 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2923 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2924 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2925 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2926 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2927 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2928 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2929 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2930 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2931 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2932 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2933 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2934 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2935 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2936 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2937 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2938 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2939 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2940 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2941 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2942 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2943 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2944 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2945 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2946 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2947 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2948 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2949 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2950 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2951 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2952 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2953 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2954 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2955 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2956 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2957 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2958 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2959 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2960 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2961 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2962 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2963 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2964 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2965 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2966 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2967 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2968 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2969 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2970 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2971 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2972 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2973 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2974 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2975 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2976 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2977 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2978 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2979 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2980 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2981 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2982 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2983 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2984 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2985 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2986 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2987 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2988 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2989 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2990 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2991 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2992 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2993 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2994 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2995 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2996 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2997 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2998 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2999 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3000 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3001 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3002 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3003 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3004 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3005 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3006 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3007 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3008 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3009 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3010 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3011 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3012 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3013 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3014 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3015 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3016 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3017 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3018 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3019 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3020 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3021 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3022 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3023 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3024 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3025 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3026 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3027 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3028 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3029 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3030 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3031 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3032 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3033 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3034 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3035 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3036 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3037 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3038 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3039 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3040 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3041 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3042 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3043 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3044 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3045 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3046 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3047 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3048 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3049 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3050 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3051 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3052 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3053 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3054 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3055 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3056 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3057 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3058 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3059 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3060 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3061 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3062 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3063 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3064 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3065 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3066 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3067 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3068 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3069 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3070 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3071 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3072 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3073 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3074 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3075 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3076 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3077 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3078 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3079 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3080 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3081 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3082 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3083 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3084 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3085 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3086 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3087 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3088 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3089 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3090 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3091 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3092 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3093 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3094 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3095 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3096 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3097 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3098 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3099 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3100 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3101 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3102 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3103 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3104 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3105 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3106 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3107 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3108 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3109 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3110 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3111 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3112 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3113 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3114 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3115 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3116 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3117 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3118 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3119 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3120 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3121 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3122 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3123 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3124 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3125 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3126 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3127 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3128 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3129 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3130 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3131 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3132 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3133 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3134 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3135 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3136 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3137 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3138 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3139 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3140 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3141 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3142 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3143 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3144 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3145 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3146 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3147 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3148 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3149 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3150 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3151 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3152 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3153 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3154 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3155 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3156 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3157 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3158 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3159 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3160 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3161 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3162 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3163 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3164 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3165 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3166 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3167 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3168 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3169 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3170 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3171 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3172 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3173 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3174 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3175 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3176 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3177 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3178 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3179 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3180 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3181 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3182 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3183 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3184 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3185 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3186 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3187 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3188 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3189 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3190 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3191 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3192 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3193 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3194 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3195 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3196 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3197 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3198 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3199 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3200 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3201 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3202 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3203 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3204 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3205 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3206 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3207 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3208 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3209 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3210 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3211 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3212 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3213 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3214 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3215 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3216 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3217 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3218 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3219 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3220 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3221 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3222 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3223 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3224 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3225 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3226 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3227 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3228 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3229 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3230 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3231 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3232 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3233 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3234 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3235 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3236 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3237 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3238 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3239 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3240 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3241 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3242 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3243 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3244 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3245 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3246 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3247 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3248 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3249 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3250 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3251 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3252 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3253 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3254 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3255 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3256 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3257 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3258 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3259 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3260 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3261 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3262 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3263 ();
 gf180mcu_fd_sc_mcu7t5v0__buf_20 input1 (.I(io_in[8]),
    .Z(net1));
 gf180mcu_fd_sc_mcu7t5v0__buf_20 input2 (.I(io_in[9]),
    .Z(net2));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output3 (.I(net3),
    .Z(io_out[16]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output4 (.I(net4),
    .Z(io_out[17]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output5 (.I(net5),
    .Z(io_out[18]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output6 (.I(net6),
    .Z(io_out[19]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output7 (.I(net7),
    .Z(io_out[20]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output8 (.I(net8),
    .Z(io_out[21]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output9 (.I(net9),
    .Z(io_out[22]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output10 (.I(net10),
    .Z(io_out[23]));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_11 (.ZN(net11));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8499__D (.I(_0003_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8501__D (.I(_0005_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8506__D (.I(_0010_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5435__A2 (.I(_0010_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5425__A2 (.I(_0010_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5409__A2 (.I(_0010_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8514__D (.I(_0018_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8528__D (.I(_0032_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8532__D (.I(_0036_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8534__D (.I(_0038_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8537__D (.I(_0041_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8542__D (.I(_0046_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8545__D (.I(_0049_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8553__D (.I(_0057_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8560__D (.I(_0064_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8561__D (.I(_0065_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8564__D (.I(_0068_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8567__D (.I(_0071_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8571__D (.I(_0075_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8572__D (.I(_0076_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8574__D (.I(_0078_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8578__D (.I(_0594_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8594__D (.I(_0610_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7841__A1 (.I(_0610_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8595__D (.I(_0611_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7831__A1 (.I(_0612_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6572__A1 (.I(_0612_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6569__A1 (.I(_0612_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3934__I (.I(_0612_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4502__A1 (.I(_0613_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3963__I (.I(_0613_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3955__I (.I(_0613_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3936__I (.I(_0613_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4572__A1 (.I(_0614_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4569__A1 (.I(_0614_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4452__A1 (.I(_0614_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3937__I (.I(_0614_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4396__A1 (.I(_0615_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4242__A1 (.I(_0615_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4239__A1 (.I(_0615_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3938__I (.I(_0615_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4441__A1 (.I(_0616_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4385__A1 (.I(_0616_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3976__I (.I(_0616_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3939__I (.I(_0616_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4380__A1 (.I(_0617_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4345__A1 (.I(_0617_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4164__A1 (.I(_0617_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3940__I (.I(_0617_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4566__A1 (.I(_0618_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4297__A1 (.I(_0618_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4152__I (.I(_0618_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3941__I (.I(_0618_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4425__A1 (.I(_0619_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4249__A1 (.I(_0619_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4234__A1 (.I(_0619_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3942__I (.I(_0619_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4698__A1 (.I(_0620_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4405__A1 (.I(_0620_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4148__I (.I(_0620_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3943__I (.I(_0620_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4256__A1 (.I(_0621_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4145__A1 (.I(_0621_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4140__A1 (.I(_0621_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3944__I (.I(_0621_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4745__A1 (.I(_0622_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4744__A1 (.I(_0622_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3954__A1 (.I(_0622_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3945__I (.I(_0622_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4752__I (.I(_0623_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4749__A1 (.I(_0623_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4192__A1 (.I(_0623_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3946__I (.I(_0623_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4787__A1 (.I(_0624_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4770__A1 (.I(_0624_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4769__A1 (.I(_0624_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3947__I (.I(_0624_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4808__A1 (.I(_0625_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4735__A1 (.I(_0625_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4602__A1 (.I(_0625_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3948__A2 (.I(_0625_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4075__I (.I(_0630_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4070__I0 (.I(_0630_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4043__C (.I(_0630_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3954__A2 (.I(_0630_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4705__A1 (.I(_0632_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4507__A1 (.I(_0632_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4388__I (.I(_0632_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3956__I (.I(_0632_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4637__A1 (.I(_0633_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4127__A1 (.I(_0633_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3987__A1 (.I(_0633_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3957__I (.I(_0633_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4703__B (.I(_0634_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4570__B (.I(_0634_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4383__A1 (.I(_0634_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3958__I (.I(_0634_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4462__A1 (.I(_0635_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4162__A1 (.I(_0635_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3982__A1 (.I(_0635_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3959__I (.I(_0635_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4686__A1 (.I(_0636_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4542__A1 (.I(_0636_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3981__A1 (.I(_0636_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3960__I (.I(_0636_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4541__A1 (.I(_0637_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4250__A1 (.I(_0637_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4137__I (.I(_0637_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3962__A1 (.I(_0637_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4195__A1 (.I(_0638_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4027__I0 (.I(_0638_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4008__I (.I(_0638_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3962__A3 (.I(_0638_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4193__A1 (.I(_0639_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4136__A1 (.I(_0639_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3971__A1 (.I(_0639_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4455__A1 (.I(_0640_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4334__A1 (.I(_0640_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3986__A1 (.I(_0640_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3964__I (.I(_0640_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4704__A1 (.I(_0641_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4337__A1 (.I(_0641_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3968__I (.I(_0641_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3965__I (.I(_0641_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4463__A1 (.I(_0642_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4393__A1 (.I(_0642_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4336__A1 (.I(_0642_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3966__I (.I(_0642_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4702__A1 (.I(_0643_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4335__C (.I(_0643_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4221__A1 (.I(_0643_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3967__A1 (.I(_0643_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4194__A1 (.I(_0644_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4135__A1 (.I(_0644_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3970__A1 (.I(_0644_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4556__A1 (.I(_0645_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4453__B (.I(_0645_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3973__I (.I(_0645_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3969__A1 (.I(_0645_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4280__A2 (.I(_0646_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4134__A1 (.I(_0646_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3970__A2 (.I(_0646_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4126__A2 (.I(_0648_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3972__A2 (.I(_0648_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4439__A1 (.I(_0650_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4309__A1 (.I(_0650_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3985__A1 (.I(_0650_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3974__I (.I(_0650_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4660__A1 (.I(_0651_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4536__A1 (.I(_0651_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4150__A1 (.I(_0651_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3975__A1 (.I(_0651_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4151__A1 (.I(_0652_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4146__A1 (.I(_0652_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3993__A1 (.I(_0652_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4555__A1 (.I(_0653_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4323__A1 (.I(_0653_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4216__I (.I(_0653_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3977__I (.I(_0653_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4537__A1 (.I(_0654_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4423__A1 (.I(_0654_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4321__A1 (.I(_0654_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3978__I (.I(_0654_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4418__A1 (.I(_0655_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4157__A1 (.I(_0655_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4155__A1 (.I(_0655_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3980__A1 (.I(_0655_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4223__A1 (.I(_0656_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4192__A2 (.I(_0656_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4145__A2 (.I(_0656_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3980__A2 (.I(_0656_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4156__A1 (.I(_0657_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4146__A2 (.I(_0657_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3993__A2 (.I(_0657_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4320__A2 (.I(_0660_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4249__A3 (.I(_0660_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4161__A1 (.I(_0660_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3991__A1 (.I(_0660_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4234__A2 (.I(_0661_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4123__A1 (.I(_0661_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4088__B (.I(_0661_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3985__A2 (.I(_0661_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4233__A1 (.I(_0662_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4172__A1 (.I(_0662_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3990__A1 (.I(_0662_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4332__A1 (.I(_0665_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4237__A1 (.I(_0665_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4171__A1 (.I(_0665_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3989__A2 (.I(_0665_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3990__A2 (.I(_0666_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4161__A2 (.I(_0667_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3991__A2 (.I(_0667_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4188__A3 (.I(_0669_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4147__A3 (.I(_0669_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3993__A3 (.I(_0669_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4125__A2 (.I(_0670_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3994__A2 (.I(_0670_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4818__A1 (.I(_0673_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4178__A2 (.I(_0673_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4119__A2 (.I(_0673_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4117__A1 (.I(_0673_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4818__A2 (.I(_0674_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4061__A1 (.I(_0674_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4028__A1 (.I(_0674_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3999__A1 (.I(_0674_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4639__A3 (.I(_0678_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4501__A1 (.I(_0678_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4022__B1 (.I(_0678_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4002__I (.I(_0678_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4640__A2 (.I(_0679_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4053__I0 (.I(_0679_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4017__A1 (.I(_0679_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4380__A2 (.I(_0680_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4044__I0 (.I(_0680_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4015__B1 (.I(_0680_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4012__A1 (.I(_0680_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4380__A3 (.I(_0682_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4031__I0 (.I(_0682_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4012__B1 (.I(_0682_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4010__I (.I(_0682_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4037__I1 (.I(_0683_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4012__B2 (.I(_0683_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4379__A1 (.I(_0687_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4279__A1 (.I(_0687_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4037__I0 (.I(_0687_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4011__A1 (.I(_0687_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4385__A2 (.I(_0691_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4049__I (.I(_0691_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4016__A2 (.I(_0691_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4015__A2 (.I(_0691_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4792__A1 (.I(_0696_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4024__A1 (.I(_0696_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4023__A1 (.I(_0696_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4022__A1 (.I(_0696_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4042__S (.I(_0702_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4036__I (.I(_0702_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4035__S (.I(_0702_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4026__I (.I(_0702_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4074__S (.I(_0703_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4063__B1 (.I(_0703_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4031__S (.I(_0703_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4027__S (.I(_0703_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4090__A2 (.I(_0708_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4079__A2 (.I(_0708_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4078__B1 (.I(_0708_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4046__A2 (.I(_0708_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4299__B2 (.I(_0709_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4140__A3 (.I(_0709_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4138__A2 (.I(_0709_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4033__I (.I(_0709_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4086__B (.I(_0710_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4073__I (.I(_0710_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4043__A1 (.I(_0710_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4040__A1 (.I(_0710_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4407__A1 (.I(_0715_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4406__A3 (.I(_0715_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4207__A2 (.I(_0715_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4039__I (.I(_0715_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4477__A2 (.I(_0716_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4408__A1 (.I(_0716_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4299__A1 (.I(_0716_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4040__B2 (.I(_0716_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4097__I1 (.I(_0721_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4079__B1 (.I(_0721_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4052__A2 (.I(_0721_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4046__C1 (.I(_0721_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4102__A1 (.I(_0727_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4055__A2 (.I(_0727_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4051__A2 (.I(_0727_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4107__A1 (.I(_0730_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4059__A2 (.I(_0730_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4055__B1 (.I(_0730_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4621__A1 (.I(_0731_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4516__A2 (.I(_0731_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4058__I (.I(_0731_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4055__B2 (.I(_0731_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4111__A1 (.I(_0740_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4067__B1 (.I(_0740_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4064__A2 (.I(_0740_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4784__A1 (.I(_0743_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4783__A1 (.I(_0743_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4112__A1 (.I(_0743_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4067__B2 (.I(_0743_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4101__I (.I(_0746_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4097__S (.I(_0746_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4089__I (.I(_0746_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4070__S (.I(_0746_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4121__A2 (.I(_0747_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4094__A1 (.I(_0747_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4184__A1 (.I(_0748_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4183__I0 (.I(_0748_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4093__B (.I(_0748_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4088__A1 (.I(_0748_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4087__A2 (.I(_0751_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4078__A2 (.I(_0751_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4076__A2 (.I(_0751_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4096__A1 (.I(_0754_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4092__A1 (.I(_0754_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4079__A1 (.I(_0754_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4078__B2 (.I(_0754_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4266__A1 (.I(_0768_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4265__I0 (.I(_0768_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4095__I (.I(_0768_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4092__C (.I(_0768_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4265__I1 (.I(_0773_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4100__A2 (.I(_0773_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4355__I1 (.I(_0774_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4105__A2 (.I(_0774_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4100__B1 (.I(_0774_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4570__C (.I(_0775_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4356__A1 (.I(_0775_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4355__I0 (.I(_0775_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4099__I (.I(_0775_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4360__A1 (.I(_0780_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4110__A2 (.I(_0780_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4106__B1 (.I(_0780_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4361__A1 (.I(_0781_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4359__A1 (.I(_0781_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4110__A1 (.I(_0781_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4106__B2 (.I(_0781_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4593__A1 (.I(_0786_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4592__A1 (.I(_0786_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4113__A1 (.I(_0786_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4110__B2 (.I(_0786_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4724__A1 (.I(_0789_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4115__B1 (.I(_0789_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4113__B1 (.I(_0789_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4187__A1 (.I(_0802_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4143__A1 (.I(_0802_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4201__A1 (.I(_0803_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4128__I (.I(_0803_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4379__A2 (.I(_0804_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4279__A2 (.I(_0804_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4194__A2 (.I(_0804_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4129__I (.I(_0804_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4504__A1 (.I(_0806_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4386__A1 (.I(_0806_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4282__A1 (.I(_0806_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4131__I (.I(_0806_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4240__I (.I(_0807_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4198__A1 (.I(_0807_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4166__A1 (.I(_0807_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4132__A1 (.I(_0807_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4287__B1 (.I(_0808_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4286__A2 (.I(_0808_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4197__A3 (.I(_0808_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4133__I (.I(_0808_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4383__B (.I(_0809_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4280__A3 (.I(_0809_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4199__A2 (.I(_0809_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4134__A2 (.I(_0809_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4191__A1 (.I(_0812_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4142__A1 (.I(_0812_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4406__A1 (.I(_0813_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4346__A1 (.I(_0813_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4207__A1 (.I(_0813_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4138__A1 (.I(_0813_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4209__A3 (.I(_0814_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4208__A2 (.I(_0814_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4139__A2 (.I(_0814_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4477__A3 (.I(_0816_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4408__A2 (.I(_0816_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4299__A2 (.I(_0816_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4141__A2 (.I(_0816_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4187__A2 (.I(_0818_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4143__A2 (.I(_0818_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4219__A1 (.I(_0820_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4192__A3 (.I(_0820_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4153__A2 (.I(_0820_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4145__A3 (.I(_0820_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4188__A2 (.I(_0822_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4147__A2 (.I(_0822_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4516__A1 (.I(_0824_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4431__A1 (.I(_0824_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4257__A1 (.I(_0824_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4149__A1 (.I(_0824_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4213__A1 (.I(_0825_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4212__A1 (.I(_0825_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4174__A1 (.I(_0825_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4420__B (.I(_0826_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4219__A2 (.I(_0826_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4151__A2 (.I(_0826_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4620__A1 (.I(_0828_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4446__A1 (.I(_0828_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4420__A1 (.I(_0828_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4153__A1 (.I(_0828_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4403__A2 (.I(_0829_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4307__A2 (.I(_0829_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4154__A2 (.I(_0829_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4215__A1 (.I(_0830_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4159__A1 (.I(_0830_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4426__A1 (.I(_0833_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4311__A2 (.I(_0833_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4158__A2 (.I(_0833_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4215__A2 (.I(_0834_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4159__A2 (.I(_0834_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4322__A3 (.I(_0838_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4319__A3 (.I(_0838_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4163__A2 (.I(_0838_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4346__A3 (.I(_0840_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4320__A3 (.I(_0840_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4165__A2 (.I(_0840_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4639__A1 (.I(_0844_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4382__A1 (.I(_0844_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4200__A1 (.I(_0844_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4169__A1 (.I(_0844_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4213__A2 (.I(_0849_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4212__A2 (.I(_0849_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4174__A3 (.I(_0849_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4189__A2 (.I(_0851_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4176__A2 (.I(_0851_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4190__A1 (.I(_0863_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4398__A1 (.I(_0871_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4392__B2 (.I(_0871_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4280__A1 (.I(_0871_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4197__A2 (.I(_0871_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4283__A1 (.I(_0875_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4201__A2 (.I(_0875_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4377__B (.I(_0877_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4281__A1 (.I(_0877_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4203__I (.I(_0877_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4378__A1 (.I(_0878_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4293__A1 (.I(_0878_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4292__A2 (.I(_0878_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4205__A1 (.I(_0878_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4278__A1 (.I(_0881_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4210__A1 (.I(_0881_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4299__B1 (.I(_0882_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4208__B (.I(_0882_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4699__A1 (.I(_0891_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4322__A1 (.I(_0891_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4306__A1 (.I(_0891_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4217__A1 (.I(_0891_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4419__A1 (.I(_0893_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4403__A1 (.I(_0893_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4307__A1 (.I(_0893_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4220__I1 (.I(_0893_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4425__A3 (.I(_0897_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4424__A1 (.I(_0897_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4311__A1 (.I(_0897_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4224__I1 (.I(_0897_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4368__A1 (.I(_0901_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4304__A1 (.I(_0901_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4301__A1 (.I(_0901_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4228__A1 (.I(_0901_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4304__B2 (.I(_0907_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4259__A1 (.I(_0907_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4454__A3 (.I(_0914_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4338__A1 (.I(_0914_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4333__A1 (.I(_0914_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4245__A2 (.I(_0914_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4454__A1 (.I(_0915_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4443__A1 (.I(_0915_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4287__A1 (.I(_0915_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4241__A1 (.I(_0915_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4330__A1 (.I(_0921_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4317__A1 (.I(_0921_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4252__A2 (.I(_0921_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4439__A3 (.I(_0922_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4320__A1 (.I(_0922_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4250__A2 (.I(_0922_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4248__I (.I(_0922_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4465__A1 (.I(_0923_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4464__A1 (.I(_0923_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4346__A2 (.I(_0923_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4251__A1 (.I(_0923_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4318__B1 (.I(_0927_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4303__A1 (.I(_0927_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4259__A2 (.I(_0927_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4551__A1 (.I(_0929_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4319__A1 (.I(_0929_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4258__A1 (.I(_0929_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4257__A2 (.I(_0929_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4446__A2 (.I(_0930_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4436__A1 (.I(_0930_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4324__A1 (.I(_0930_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4256__A2 (.I(_0930_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4318__B2 (.I(_0933_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4303__A2 (.I(_0933_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4259__A3 (.I(_0933_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4637__A2 (.I(_0958_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4505__A1 (.I(_0958_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4396__A2 (.I(_0958_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4285__I (.I(_0958_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4376__A2 (.I(_0965_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4375__A2 (.I(_0965_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4296__A1 (.I(_0965_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4376__A1 (.I(_0966_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4295__A1 (.I(_0966_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4294__A2 (.I(_0966_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4375__A1 (.I(_0968_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4295__A2 (.I(_0968_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4374__A2 (.I(_0974_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4367__A2 (.I(_0974_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4301__A3 (.I(_0974_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4542__C (.I(_0980_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4419__A2 (.I(_0980_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4403__A3 (.I(_0980_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4308__A1 (.I(_0980_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4416__A1 (.I(_0982_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4313__A1 (.I(_0982_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4537__C (.I(_0983_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4310__I (.I(_0983_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4482__A1 (.I(_0988_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4414__B2 (.I(_0988_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4411__A1 (.I(_0988_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4316__A1 (.I(_0988_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4414__A1 (.I(_0992_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4349__A1 (.I(_0992_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4437__A1 (.I(_0993_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4327__A1 (.I(_0993_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4326__A1 (.I(_0993_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4681__A2 (.I(_0995_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4554__A2 (.I(_0995_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4436__A2 (.I(_0995_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4324__A2 (.I(_0995_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4689__A3 (.I(_0997_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4440__A2 (.I(_0997_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4436__B2 (.I(_0997_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4324__B2 (.I(_0997_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4437__A2 (.I(_0999_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4327__A2 (.I(_0999_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4326__A2 (.I(_0999_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4413__A1 (.I(_1002_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4412__A1 (.I(_1002_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4349__A2 (.I(_1002_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4330__B (.I(_1003_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4449__A1 (.I(_1007_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4342__A1 (.I(_1007_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4449__A2 (.I(_1015_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4342__A2 (.I(_1015_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4580__B2 (.I(_1017_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4462__A2 (.I(_1017_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4345__A2 (.I(_1017_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4344__I (.I(_1017_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4464__A2 (.I(_1019_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4439__A4 (.I(_1019_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4347__I1 (.I(_1019_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4413__A2 (.I(_1022_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4412__A2 (.I(_1022_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4349__A3 (.I(_1022_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4372__A2 (.I(_1024_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4364__A2 (.I(_1024_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4351__A3 (.I(_1024_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4723__A1 (.I(_1031_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4594__A1 (.I(_1031_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4476__A1 (.I(_1031_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4475__A1 (.I(_1031_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4494__A1 (.I(_1052_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4402__A1 (.I(_1052_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4645__A1 (.I(_1061_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4640__B (.I(_1061_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4579__I (.I(_1061_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4392__A1 (.I(_1061_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4637__A3 (.I(_1062_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4504__A2 (.I(_1062_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4393__A3 (.I(_1062_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4390__I (.I(_1062_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4644__A1 (.I(_1063_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4642__A1 (.I(_1063_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4396__A3 (.I(_1063_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4392__A2 (.I(_1063_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4507__B1 (.I(_1064_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4499__A2 (.I(_1064_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4398__A2 (.I(_1064_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4392__B1 (.I(_1064_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4496__C (.I(_1072_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4495__A2 (.I(_1072_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4400__A2 (.I(_1072_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4494__A2 (.I(_1074_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4402__A2 (.I(_1074_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4492__A1 (.I(_1075_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4491__A1 (.I(_1075_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4404__A2 (.I(_1075_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4492__A2 (.I(_1076_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4491__A2 (.I(_1076_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4404__A3 (.I(_1076_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4490__A2 (.I(_1082_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4410__A3 (.I(_1082_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4416__A2 (.I(_1088_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4661__A1 (.I(_1090_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4660__A3 (.I(_1090_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4513__I (.I(_1090_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4418__A2 (.I(_1090_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4543__A2 (.I(_1091_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4422__A1 (.I(_1091_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4628__A2 (.I(_1093_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4627__A2 (.I(_1093_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4514__A2 (.I(_1093_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4421__A2 (.I(_1093_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4533__B2 (.I(_1095_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4429__A1 (.I(_1095_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4538__A2 (.I(_1096_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4428__A1 (.I(_1096_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4427__A1 (.I(_1097_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4426__A2 (.I(_1097_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4528__A1 (.I(_1108_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4527__A1 (.I(_1108_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4468__A2 (.I(_1108_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4438__A1 (.I(_1109_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4551__A2 (.I(_1113_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4444__A2 (.I(_1113_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4557__A2 (.I(_1114_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4556__B1 (.I(_1114_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4446__A4 (.I(_1114_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4442__A2 (.I(_1114_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4549__A1 (.I(_1122_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4548__A1 (.I(_1122_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4467__A2 (.I(_1122_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4565__A1 (.I(_1124_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4460__A1 (.I(_1124_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4704__A3 (.I(_1125_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4573__A1 (.I(_1125_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4459__A1 (.I(_1125_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4565__A2 (.I(_1132_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4460__A2 (.I(_1132_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4769__A2 (.I(_1134_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4697__A1 (.I(_1134_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4696__A1 (.I(_1134_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4462__A3 (.I(_1134_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4581__A3 (.I(_1136_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4580__B1 (.I(_1136_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4555__A4 (.I(_1136_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4464__B (.I(_1136_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4528__A2 (.I(_1140_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4527__A2 (.I(_1140_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4468__A3 (.I(_1140_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4485__A2 (.I(_1141_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4484__A2 (.I(_1141_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4469__A2 (.I(_1141_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4601__A1 (.I(_1149_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4588__A1 (.I(_1149_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4607__A1 (.I(_1162_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4525__A2 (.I(_1162_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4630__A1 (.I(_1169_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4512__A1 (.I(_1169_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4799__A2 (.I(_1176_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4798__A2 (.I(_1176_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4505__A2 (.I(_1176_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4630__A2 (.I(_1183_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4512__A2 (.I(_1183_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4754__A1 (.I(_1185_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4628__A1 (.I(_1185_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4627__A1 (.I(_1185_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4514__A1 (.I(_1185_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4613__A2 (.I(_1187_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4612__A2 (.I(_1187_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4524__A2 (.I(_1187_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4614__A2 (.I(_1195_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4524__A3 (.I(_1195_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4664__A1 (.I(_1202_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4531__I (.I(_1202_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4751__A1 (.I(_1203_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4668__A1 (.I(_1203_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4534__A1 (.I(_1203_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4533__A1 (.I(_1203_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4615__A1 (.I(_1205_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4547__A1 (.I(_1205_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4657__A1 (.I(_1206_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4535__I (.I(_1206_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4751__A3 (.I(_1208_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4658__A1 (.I(_1208_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4540__A1 (.I(_1208_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4738__A2 (.I(_1209_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4671__A2 (.I(_1209_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4539__A1 (.I(_1209_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4657__A2 (.I(_1212_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4546__A2 (.I(_1212_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4755__B1 (.I(_1213_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4545__A1 (.I(_1213_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4632__A2 (.I(_1214_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4544__A1 (.I(_1214_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4658__B2 (.I(_1217_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4546__A3 (.I(_1217_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4680__A1 (.I(_1227_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4559__A1 (.I(_1227_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4680__A2 (.I(_1230_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4559__A2 (.I(_1230_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4788__A1 (.I(_1234_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4674__A1 (.I(_1234_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4564__A1 (.I(_1234_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4694__A1 (.I(_1249_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4582__A1 (.I(_1249_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4763__A1 (.I(_1251_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4666__A1 (.I(_1251_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4662__B (.I(_1251_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4580__A1 (.I(_1251_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4610__A2 (.I(_1257_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4609__A2 (.I(_1257_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4586__A3 (.I(_1257_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4604__A2 (.I(_1258_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4603__A2 (.I(_1258_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4587__A3 (.I(_1258_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4594__A2 (.I(_1262_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4726__B2 (.I(_1273_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4719__A1 (.I(_1273_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4761__A1 (.I(_1285_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4653__A1 (.I(_1285_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4736__A1 (.I(_1293_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4626__A1 (.I(_1293_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4777__A1 (.I(_1297_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4651__A1 (.I(_1297_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4776__A1 (.I(_1300_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4775__A1 (.I(_1300_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4651__A2 (.I(_1300_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4776__A2 (.I(_1321_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4775__A2 (.I(_1321_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4651__A3 (.I(_1321_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4760__A2 (.I(_1322_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4652__A2 (.I(_1322_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4739__A1 (.I(_1334_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4673__A1 (.I(_1334_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4665__A2 (.I(_1335_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4741__I (.I(_1338_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4738__A1 (.I(_1338_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4671__A1 (.I(_1338_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4668__A2 (.I(_1338_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4670__A1 (.I(_1339_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4669__A2 (.I(_1339_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4751__B (.I(_1340_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4670__B (.I(_1340_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4672__S (.I(_1342_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4788__A2 (.I(_1344_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4674__A2 (.I(_1344_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4771__A1 (.I(_1354_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4763__A2 (.I(_1354_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4689__A2 (.I(_1354_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4684__A2 (.I(_1354_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4694__B (.I(_1364_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4769__A4 (.I(_1366_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4733__A2 (.I(_1366_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4697__A3 (.I(_1366_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4696__B (.I(_1366_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4809__A1 (.I(_1372_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4710__A1 (.I(_1372_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4746__A2 (.I(_1376_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4706__A2 (.I(_1376_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4809__A2 (.I(_1380_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4710__A2 (.I(_1380_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4726__A2 (.I(_1388_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4718__A2 (.I(_1388_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4735__A2 (.I(_1404_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4740__A1 (.I(_1407_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4742__A1 (.I(_1411_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4743__A2 (.I(_1412_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4793__A1 (.I(_1422_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4767__B (.I(_1422_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4766__A1 (.I(_1422_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4757__A1 (.I(_1422_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4794__A1 (.I(_1423_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4755__A2 (.I(_1423_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4754__A2 (.I(_1423_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4758__A2 (.I(_1427_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4762__A2 (.I(_1429_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4774__A2 (.I(_1438_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4803__A1 (.I(_1444_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4782__A2 (.I(_1451_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4787__A2 (.I(_1456_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4802__A2 (.I(_1457_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4801__A1 (.I(_1459_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4793__A2 (.I(_1462_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4801__A2 (.I(_1463_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4800__A3 (.I(_1469_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4804__A3 (.I(_1473_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4814__A2 (.I(_1483_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6390__S0 (.I(_1489_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5420__I (.I(_1489_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4956__I (.I(_1489_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4821__I (.I(_1489_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6272__C (.I(_1490_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5788__A1 (.I(_1490_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5195__C (.I(_1490_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4822__I (.I(_1490_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6548__A1 (.I(_1491_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6509__A1 (.I(_1491_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5790__A1 (.I(_1491_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4961__A1 (.I(_1491_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6292__I (.I(_1493_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5634__I (.I(_1493_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5578__I (.I(_1493_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4828__A1 (.I(_1493_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6068__B (.I(_1495_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5457__I (.I(_1495_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4830__I (.I(_1495_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4827__A2 (.I(_1495_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6125__A2 (.I(_1497_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6084__A2 (.I(_1497_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4829__I (.I(_1497_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5872__C (.I(_1498_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5840__C (.I(_1498_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5747__C (.I(_1498_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4961__A2 (.I(_1498_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5731__A2 (.I(_1499_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5089__I (.I(_1499_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4950__I (.I(_1499_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4837__A1 (.I(_1499_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5403__I (.I(_1501_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4957__A1 (.I(_1501_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4860__A1 (.I(_1501_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4836__A1 (.I(_1501_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5249__I (.I(_1503_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5145__I (.I(_1503_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4872__A2 (.I(_1503_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4835__A2 (.I(_1503_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4892__A2 (.I(_1504_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4880__I (.I(_1504_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4855__A1 (.I(_1504_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4836__A2 (.I(_1504_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6120__A1 (.I(_1505_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6117__A2 (.I(_1505_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4837__A2 (.I(_1505_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5319__B (.I(_1508_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5110__C (.I(_1508_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5088__A1 (.I(_1508_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4878__A1 (.I(_1508_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5304__I (.I(_1509_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4981__S (.I(_1509_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4940__I (.I(_1509_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4841__I (.I(_1509_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5477__S (.I(_1510_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5142__S (.I(_1510_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5140__S (.I(_1510_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4842__S (.I(_1510_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5278__I (.I(_1514_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5007__I (.I(_1514_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4871__S (.I(_1514_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4846__I (.I(_1514_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5985__S (.I(_1515_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5743__S (.I(_1515_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5306__S (.I(_1515_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4847__S (.I(_1515_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6123__A2 (.I(_1516_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4863__I2 (.I(_1516_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5794__I (.I(_1517_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5698__I (.I(_1517_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5147__I (.I(_1517_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4849__I (.I(_1517_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5115__I (.I(_1518_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5079__I (.I(_1518_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5017__I (.I(_1518_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4850__I (.I(_1518_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5828__I (.I(_1519_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5076__S (.I(_1519_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4988__S (.I(_1519_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4851__S (.I(_1519_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6123__B1 (.I(_1520_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4863__I3 (.I(_1520_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5447__I (.I(_1522_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5398__I (.I(_1522_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5022__I (.I(_1522_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4854__A1 (.I(_1522_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5084__I (.I(_1524_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5075__I (.I(_1524_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4856__I (.I(_1524_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4995__I (.I(_1525_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4933__I (.I(_1525_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4895__I (.I(_1525_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4857__I (.I(_1525_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5519__I (.I(_1527_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5318__S0 (.I(_1527_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5129__S0 (.I(_1527_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4863__S0 (.I(_1527_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4902__A1 (.I(_1528_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4868__I (.I(_1528_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4860__A2 (.I(_1528_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4973__I (.I(_1529_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4861__I (.I(_1529_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5217__I (.I(_1530_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5156__I (.I(_1530_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5128__I (.I(_1530_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4862__I (.I(_1530_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5167__B (.I(_1531_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4994__B (.I(_1531_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4876__B1 (.I(_1531_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4863__S1 (.I(_1531_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4878__A2 (.I(_1532_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5945__A1 (.I(_1533_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5748__A2 (.I(_1533_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5545__I (.I(_1533_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4878__B (.I(_1533_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6064__B (.I(_1535_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5851__I (.I(_1535_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5451__I (.I(_1535_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4867__I (.I(_1535_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6431__A1 (.I(_1536_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5959__B (.I(_1536_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4890__A2 (.I(_1536_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4877__A1 (.I(_1536_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6288__I (.I(_1537_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5062__I (.I(_1537_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4886__A2 (.I(_1537_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4869__I (.I(_1537_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6386__A2 (.I(_1538_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6135__I (.I(_1538_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5561__I (.I(_1538_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4870__I (.I(_1538_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6114__A2 (.I(_1539_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5552__A2 (.I(_1539_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4959__A1 (.I(_1539_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4876__A2 (.I(_1539_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6096__A2 (.I(_1541_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4902__A2 (.I(_1541_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4873__I (.I(_1541_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6089__A2 (.I(_1542_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5748__A1 (.I(_1542_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5562__I (.I(_1542_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4874__I (.I(_1542_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6289__I (.I(_1543_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5516__I (.I(_1543_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5143__I (.I(_1543_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4875__S (.I(_1543_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5777__A2 (.I(_1548_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5571__I (.I(_1548_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5443__I (.I(_1548_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4881__A1 (.I(_1548_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5589__I (.I(_1549_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5583__I (.I(_1549_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5431__I (.I(_1549_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4881__A2 (.I(_1549_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5319__A1 (.I(_1551_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5284__A1 (.I(_1551_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4890__C (.I(_1551_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4883__I (.I(_1551_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5247__A1 (.I(_1552_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5196__A1 (.I(_1552_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5003__A1 (.I(_1552_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4891__A2 (.I(_1552_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5729__A2 (.I(_1553_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5404__A2 (.I(_1553_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4957__A2 (.I(_1553_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4887__A1 (.I(_1553_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5770__A2 (.I(_1554_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5452__A2 (.I(_1554_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4892__A1 (.I(_1554_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4886__A1 (.I(_1554_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6204__B2 (.I(_1555_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6164__A1 (.I(_1555_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4887__A2 (.I(_1555_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5197__I (.I(_1557_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5155__A1 (.I(_1557_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5144__C (.I(_1557_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4889__I (.I(_1557_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5131__C (.I(_1558_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5029__B (.I(_1558_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4923__B (.I(_1558_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4890__B2 (.I(_1558_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4961__A3 (.I(_1560_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4983__I (.I(_1561_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4945__I (.I(_1561_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4921__I (.I(_1561_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4893__I (.I(_1561_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5081__B (.I(_1562_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5073__B (.I(_1562_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5032__I (.I(_1562_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4894__I (.I(_1562_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5275__C (.I(_1563_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5107__A1 (.I(_1563_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4948__A1 (.I(_1563_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4908__A1 (.I(_1563_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6290__I (.I(_1564_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6136__I (.I(_1564_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4915__I (.I(_1564_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4896__I (.I(_1564_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6385__A1 (.I(_1565_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5096__S (.I(_1565_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4982__A1 (.I(_1565_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4897__I (.I(_1565_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6320__A1 (.I(_1566_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6204__A1 (.I(_1566_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6164__B2 (.I(_1566_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4901__A1 (.I(_1566_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5116__I (.I(_1567_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5039__I (.I(_1567_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4943__I (.I(_1567_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4899__I (.I(_1567_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5317__S (.I(_1568_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5314__S (.I(_1568_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4935__S (.I(_1568_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4900__S (.I(_1568_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5027__I (.I(_1571_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4903__I (.I(_1571_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6145__I (.I(_1573_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5276__I (.I(_1573_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5036__I (.I(_1573_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4905__I (.I(_1573_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6257__I (.I(_1574_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5599__A1 (.I(_1574_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5152__A1 (.I(_1574_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4906__I (.I(_1574_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6120__B2 (.I(_1575_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6117__B1 (.I(_1575_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4914__A1 (.I(_1575_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4907__A2 (.I(_1575_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5179__I (.I(_1578_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5046__I (.I(_1578_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4917__I (.I(_1578_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4910__I (.I(_1578_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5289__I (.I(_1579_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5112__I (.I(_1579_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5024__I (.I(_1579_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4911__I (.I(_1579_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5353__S (.I(_1580_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5257__S (.I(_1580_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5212__I (.I(_1580_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4912__I (.I(_1580_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5764__S (.I(_1581_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5703__I (.I(_1581_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5166__S (.I(_1581_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4913__S (.I(_1581_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6102__A2 (.I(_1582_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4914__A2 (.I(_1582_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6364__A1 (.I(_1585_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6226__A1 (.I(_1585_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6179__A1 (.I(_1585_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4922__A1 (.I(_1585_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5758__I (.I(_1588_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5370__S (.I(_1588_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5224__S (.I(_1588_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4920__S (.I(_1588_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6103__A2 (.I(_1589_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4922__A2 (.I(_1589_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5383__S1 (.I(_1590_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5367__S1 (.I(_1590_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5343__S1 (.I(_1590_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4922__B (.I(_1590_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5596__I (.I(_1594_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5018__I (.I(_1594_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4968__I (.I(_1594_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4928__A1 (.I(_1594_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5770__A1 (.I(_1595_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5750__A1 (.I(_1595_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5410__I (.I(_1595_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4927__A1 (.I(_1595_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5303__A2 (.I(_1599_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5297__A2 (.I(_1599_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5266__A2 (.I(_1599_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4949__B (.I(_1599_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5590__I (.I(_1600_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5082__I (.I(_1600_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4971__I (.I(_1600_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4932__I (.I(_1600_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5574__I (.I(_1601_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5141__A2 (.I(_1601_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5066__A2 (.I(_1601_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4936__A2 (.I(_1601_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6319__A1 (.I(_1603_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5106__A1 (.I(_1603_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4946__A1 (.I(_1603_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4936__B1 (.I(_1603_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4948__A2 (.I(_1605_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5591__I (.I(_1606_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5070__I (.I(_1606_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4976__I (.I(_1606_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4938__I (.I(_1606_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5382__I (.I(_1607_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5216__I (.I(_1607_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5097__I (.I(_1607_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4939__I (.I(_1607_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6345__A1 (.I(_1608_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5165__A1 (.I(_1608_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4992__A1 (.I(_1608_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4942__A1 (.I(_1608_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5900__I (.I(_1609_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5657__I (.I(_1609_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5326__S (.I(_1609_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4941__S (.I(_1609_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6088__A2 (.I(_1610_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4942__A2 (.I(_1610_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6049__A1 (.I(_1612_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5800__I (.I(_1612_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5286__S (.I(_1612_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4944__S (.I(_1612_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6092__A2 (.I(_1613_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4946__A2 (.I(_1613_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5184__A1 (.I(_1614_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5165__B (.I(_1614_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4992__B (.I(_1614_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4946__B (.I(_1614_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5087__C (.I(_1616_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4999__C (.I(_1616_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4965__I (.I(_1616_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4948__C (.I(_1616_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4955__A1 (.I(_1618_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6084__B2 (.I(_1620_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5989__A1 (.I(_1620_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4966__A1 (.I(_1620_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4954__A1 (.I(_1620_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5375__B (.I(_1621_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5199__A2 (.I(_1621_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5195__A1 (.I(_1621_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4954__B1 (.I(_1621_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5312__A1 (.I(_1622_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5296__A1 (.I(_1622_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5000__B (.I(_1622_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4954__C (.I(_1622_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4961__B1 (.I(_1624_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6141__C (.I(_1625_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6125__C (.I(_1625_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5199__B (.I(_1625_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4960__A1 (.I(_1625_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6250__A2 (.I(_1627_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5965__A1 (.I(_1627_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5135__A2 (.I(_1627_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4959__A2 (.I(_1627_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5234__A2 (.I(_1628_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4963__I (.I(_1628_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4960__A2 (.I(_1628_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5395__C (.I(_1629_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5358__C (.I(_1629_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5263__C (.I(_1629_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4961__B2 (.I(_1629_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5568__B (.I(_1631_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5299__A1 (.I(_1631_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5203__A1 (.I(_1631_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5060__A1 (.I(_1631_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7250__I0 (.I(_1632_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5834__I1 (.I(_1632_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5550__B1 (.I(_1632_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4966__A2 (.I(_1632_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5336__B (.I(_1633_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5298__A1 (.I(_1633_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5232__B (.I(_1633_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4966__B1 (.I(_1633_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6344__A1 (.I(_1635_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6337__A1 (.I(_1635_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6335__A1 (.I(_1635_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4970__A1 (.I(_1635_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5801__I (.I(_1636_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5064__S (.I(_1636_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4997__S (.I(_1636_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4969__S (.I(_1636_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6146__A2 (.I(_1637_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4970__A2 (.I(_1637_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4986__A1 (.I(_1638_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5618__B1 (.I(_1639_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5556__I (.I(_1639_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4993__I (.I(_1639_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4972__I (.I(_1639_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6148__A1 (.I(_1640_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6108__A1 (.I(_1640_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5543__B1 (.I(_1640_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4975__A2 (.I(_1640_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5374__S1 (.I(_1642_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5259__C (.I(_1642_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5193__A1 (.I(_1642_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4975__B (.I(_1642_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6171__A1 (.I(_1645_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5274__A1 (.I(_1645_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5144__A2 (.I(_1645_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4984__A1 (.I(_1645_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5210__I (.I(_1646_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5047__I (.I(_1646_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4990__I (.I(_1646_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4979__I (.I(_1646_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5186__A1 (.I(_1647_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5181__A1 (.I(_1647_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5072__S (.I(_1647_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4980__S (.I(_1647_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6150__A2 (.I(_1648_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4984__A2 (.I(_1648_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6151__A2 (.I(_1649_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4982__A2 (.I(_1649_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5106__B (.I(_1651_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5051__B (.I(_1651_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5028__S1 (.I(_1651_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4984__C (.I(_1651_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5262__I (.I(_1653_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5219__I (.I(_1653_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5157__A1 (.I(_1653_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4986__C (.I(_1653_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6373__A1 (.I(_1655_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6305__A1 (.I(_1655_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6262__A1 (.I(_1655_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4989__A1 (.I(_1655_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6155__A2 (.I(_1656_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4989__A2 (.I(_1656_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5773__I (.I(_1658_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5190__A1 (.I(_1658_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5068__S (.I(_1658_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4991__S (.I(_1658_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6154__A2 (.I(_1659_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4992__A2 (.I(_1659_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6259__I (.I(_1663_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5168__I (.I(_1663_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5160__I (.I(_1663_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4996__I (.I(_1663_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6304__A1 (.I(_1664_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6246__B1 (.I(_1664_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5566__A1 (.I(_1664_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4998__A1 (.I(_1664_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5000__A2 (.I(_1667_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5003__B (.I(_1668_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5200__I (.I(_1669_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5137__A1 (.I(_1669_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5132__I (.I(_1669_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5002__I (.I(_1669_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6175__A1 (.I(_1670_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6028__A1 (.I(_1670_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5135__B2 (.I(_1670_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5003__C (.I(_1670_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5377__A2 (.I(_1673_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5323__A2 (.I(_1673_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5206__A2 (.I(_1673_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5030__A2 (.I(_1673_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6563__A2 (.I(_1674_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5260__B (.I(_1674_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5054__A1 (.I(_1674_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5029__A1 (.I(_1674_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6068__A1 (.I(_1676_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5033__I (.I(_1676_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5013__I (.I(_1676_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5009__I (.I(_1676_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5735__I (.I(_1677_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5506__A1 (.I(_1677_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5494__A1 (.I(_1677_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5011__A1 (.I(_1677_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6171__A2 (.I(_1680_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5028__I0 (.I(_1680_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6001__I (.I(_1681_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5733__I (.I(_1681_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5316__S (.I(_1681_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5015__A1 (.I(_1681_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6172__A2 (.I(_1684_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5028__I1 (.I(_1684_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6016__A1 (.I(_1685_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5968__I (.I(_1685_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5161__S (.I(_1685_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5021__A1 (.I(_1685_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5986__S (.I(_1686_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5664__I (.I(_1686_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5497__A1 (.I(_1686_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5020__A1 (.I(_1686_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6111__I (.I(_1691_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5717__I (.I(_1691_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5684__I (.I(_1691_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5026__A1 (.I(_1691_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5671__I (.I(_1692_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5269__I (.I(_1692_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5035__S (.I(_1692_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5025__A1 (.I(_1692_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5311__S0 (.I(_1695_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5267__I (.I(_1695_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5136__I (.I(_1695_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5028__S0 (.I(_1695_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5029__A2 (.I(_1696_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5030__B (.I(_1697_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5338__A2 (.I(_1699_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5237__A2 (.I(_1699_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5202__C (.I(_1699_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5055__A2 (.I(_1699_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5386__A1 (.I(_1700_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5348__A1 (.I(_1700_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5252__A1 (.I(_1700_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5052__A1 (.I(_1700_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5424__I (.I(_1701_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5102__I (.I(_1701_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5085__S (.I(_1701_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5034__S (.I(_1701_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6164__A2 (.I(_1702_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5037__I0 (.I(_1702_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6164__B1 (.I(_1703_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5037__I1 (.I(_1703_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5391__A1 (.I(_1704_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5354__A1 (.I(_1704_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5258__A1 (.I(_1704_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5037__S (.I(_1704_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6211__A1 (.I(_1706_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6205__A1 (.I(_1706_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6165__A1 (.I(_1706_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5044__A1 (.I(_1706_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6115__S (.I(_1707_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5889__I (.I(_1707_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5100__A1 (.I(_1707_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5043__A1 (.I(_1707_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5331__S (.I(_1708_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5104__A1 (.I(_1708_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5099__A1 (.I(_1708_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5042__A1 (.I(_1708_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6166__A2 (.I(_1711_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5044__A2 (.I(_1711_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6350__S (.I(_1713_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6123__B2 (.I(_1713_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5528__I (.I(_1713_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5051__A1 (.I(_1713_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5739__S0 (.I(_1714_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5719__I (.I(_1714_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5122__A1 (.I(_1714_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5050__A1 (.I(_1714_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5513__A1 (.I(_1715_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5126__A1 (.I(_1715_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5121__A1 (.I(_1715_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5049__A1 (.I(_1715_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5201__B2 (.I(_1721_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5194__A1 (.I(_1721_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5091__B1 (.I(_1721_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5054__B (.I(_1721_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5055__B (.I(_1722_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6394__I (.I(_1724_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5405__A1 (.I(_1724_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5300__I (.I(_1724_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5057__I (.I(_1724_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6352__C (.I(_1725_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5429__I (.I(_1725_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5414__I (.I(_1725_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5058__I (.I(_1725_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6127__A1 (.I(_1726_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6078__B (.I(_1726_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5913__I (.I(_1726_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5059__B (.I(_1726_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5061__I (.I(_1728_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6228__A2 (.I(_1729_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6071__B (.I(_1729_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5533__A2 (.I(_1729_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5135__A1 (.I(_1729_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6206__A1 (.I(_1730_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6166__A1 (.I(_1730_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5141__B1 (.I(_1730_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5065__A1 (.I(_1730_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6190__A2 (.I(_1731_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5065__A2 (.I(_1731_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6222__A1 (.I(_1734_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6212__A1 (.I(_1734_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6172__A1 (.I(_1734_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5069__A1 (.I(_1734_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6193__A2 (.I(_1735_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5069__A2 (.I(_1735_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6263__I (.I(_1737_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6106__I (.I(_1737_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5617__A1 (.I(_1737_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5071__I (.I(_1737_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6370__S (.I(_1738_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6342__S (.I(_1738_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6310__S (.I(_1738_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5073__A1 (.I(_1738_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6192__A2 (.I(_1739_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5073__A2 (.I(_1739_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6270__S (.I(_1742_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6192__A1 (.I(_1742_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6150__A1 (.I(_1742_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5077__A1 (.I(_1742_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6197__A2 (.I(_1743_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5077__A2 (.I(_1743_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5295__S0 (.I(_1745_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5188__A1 (.I(_1745_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5177__A1 (.I(_1745_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5081__A1 (.I(_1745_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5616__A1 (.I(_1746_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5095__S (.I(_1746_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5094__S (.I(_1746_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5080__S (.I(_1746_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6196__A2 (.I(_1747_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5081__A2 (.I(_1747_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5614__B1 (.I(_1749_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5607__B1 (.I(_1749_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5600__B1 (.I(_1749_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5083__A2 (.I(_1749_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6196__A1 (.I(_1751_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6154__A1 (.I(_1751_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5231__S0 (.I(_1751_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5086__A1 (.I(_1751_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5093__I0 (.I(_1755_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6081__I (.I(_1756_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5899__S1 (.I(_1756_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5739__S1 (.I(_1756_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5090__I (.I(_1756_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6557__B (.I(_1757_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6007__I (.I(_1757_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5201__A1 (.I(_1757_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5091__A1 (.I(_1757_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5313__A2 (.I(_1759_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5131__A1 (.I(_1759_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5110__A1 (.I(_1759_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5093__S (.I(_1759_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5135__B1 (.I(_1760_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6204__A2 (.I(_1761_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5096__I0 (.I(_1761_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6204__B1 (.I(_1762_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5096__I1 (.I(_1762_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6103__A1 (.I(_1764_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6092__A1 (.I(_1764_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5167__A1 (.I(_1764_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5101__A1 (.I(_1764_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6206__A2 (.I(_1767_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5101__A2 (.I(_1767_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6055__S (.I(_1769_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5782__S (.I(_1769_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5309__A1 (.I(_1769_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5105__A1 (.I(_1769_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7294__A1 (.I(_1770_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6452__A2 (.I(_1770_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5104__A2 (.I(_1770_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6205__A2 (.I(_1772_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5106__A2 (.I(_1772_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5110__A2 (.I(_1774_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5393__B (.I(_1775_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5356__B (.I(_1775_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5130__A2 (.I(_1775_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5109__A2 (.I(_1775_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6000__I (.I(_1778_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5948__A1 (.I(_1778_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5498__A1 (.I(_1778_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5114__A1 (.I(_1778_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5651__I (.I(_1779_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5510__I (.I(_1779_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5253__I (.I(_1779_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5113__A1 (.I(_1779_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6209__A2 (.I(_1781_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5129__I0 (.I(_1781_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6119__S (.I(_1782_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5541__A1 (.I(_1782_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5530__I (.I(_1782_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5119__A1 (.I(_1782_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5919__I (.I(_1783_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5294__S (.I(_1783_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5273__S (.I(_1783_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5118__A1 (.I(_1783_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6210__A2 (.I(_1786_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5129__I1 (.I(_1786_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7600__A1 (.I(_1787_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5843__A2 (.I(_1787_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5121__A2 (.I(_1787_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6212__A2 (.I(_1789_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5129__I2 (.I(_1789_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5549__I (.I(_1790_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5227__I (.I(_1790_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5214__I (.I(_1790_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5124__I (.I(_1790_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5779__S (.I(_1791_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5504__A1 (.I(_1791_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5491__A1 (.I(_1791_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5127__A1 (.I(_1791_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6211__A2 (.I(_1794_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5129__I3 (.I(_1794_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6123__A1 (.I(_1795_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5318__S1 (.I(_1795_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5311__S1 (.I(_1795_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5129__S1 (.I(_1795_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5131__A2 (.I(_1796_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5486__A1 (.I(_1799_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5233__I (.I(_1799_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5138__I (.I(_1799_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5133__I (.I(_1799_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6215__A1 (.I(_1800_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5910__C (.I(_1800_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5588__A1 (.I(_1800_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5134__B (.I(_1800_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5135__C (.I(_1801_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6233__A1 (.I(_1802_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6083__A1 (.I(_1802_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5427__A1 (.I(_1802_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5204__A1 (.I(_1802_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5655__A2 (.I(_1803_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5480__A1 (.I(_1803_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5464__I (.I(_1803_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5204__A2 (.I(_1803_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5870__B (.I(_1804_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5838__B (.I(_1804_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5544__I (.I(_1804_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5159__A1 (.I(_1804_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6113__B (.I(_1805_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5283__A1 (.I(_1805_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5246__S1 (.I(_1805_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5158__A1 (.I(_1805_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5141__B2 (.I(_1806_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5144__B1 (.I(_1808_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6130__B1 (.I(_1809_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6114__B1 (.I(_1809_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5552__B1 (.I(_1809_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5144__B2 (.I(_1809_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5637__I (.I(_1811_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5597__I (.I(_1811_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5592__I (.I(_1811_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5146__I (.I(_1811_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5729__A1 (.I(_1812_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5521__I (.I(_1812_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5468__I (.I(_1812_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5149__S0 (.I(_1812_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5852__I (.I(_1814_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5378__S (.I(_1814_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5339__S (.I(_1814_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5149__S1 (.I(_1814_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5157__A2 (.I(_1815_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5287__I (.I(_1816_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5163__I (.I(_1816_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5153__S (.I(_1816_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5151__S (.I(_1816_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6224__A2 (.I(_1817_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5152__A2 (.I(_1817_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6222__A2 (.I(_1819_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5154__A2 (.I(_1819_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5155__A3 (.I(_1820_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5392__C (.I(_1822_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5355__C (.I(_1822_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5295__S1 (.I(_1822_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5157__C (.I(_1822_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5196__A2 (.I(_1825_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6313__A1 (.I(_1826_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6277__A1 (.I(_1826_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5282__A1 (.I(_1826_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5162__A1 (.I(_1826_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6235__A2 (.I(_1827_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5162__A2 (.I(_1827_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5385__S0 (.I(_1829_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5347__S0 (.I(_1829_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5251__S0 (.I(_1829_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5164__S (.I(_1829_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6234__A2 (.I(_1830_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5165__A2 (.I(_1830_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6233__A2 (.I(_1832_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5167__A2 (.I(_1832_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6367__A1 (.I(_1834_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6185__A1 (.I(_1834_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5259__A1 (.I(_1834_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5172__A1 (.I(_1834_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5340__S (.I(_1836_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5240__S (.I(_1836_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5191__A1 (.I(_1836_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5171__S (.I(_1836_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6231__A2 (.I(_1837_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5172__A2 (.I(_1837_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6064__A1 (.I(_1840_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5760__I (.I(_1840_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5631__I (.I(_1840_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5176__A1 (.I(_1840_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5374__S0 (.I(_1844_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5335__S0 (.I(_1844_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5192__A1 (.I(_1844_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5183__A1 (.I(_1844_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5625__I (.I(_1845_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5481__S (.I(_1845_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5187__A1 (.I(_1845_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5182__A1 (.I(_1845_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5894__A2 (.I(_1846_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5181__A2 (.I(_1846_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6237__A2 (.I(_1848_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5183__A2 (.I(_1848_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6240__A2 (.I(_1853_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5188__A2 (.I(_1853_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7296__A1 (.I(_1855_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6479__A2 (.I(_1855_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5190__A2 (.I(_1855_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5196__A3 (.I(_1861_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5368__B (.I(_1863_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5329__B (.I(_1863_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5312__B (.I(_1863_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5198__A2 (.I(_1863_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6382__C (.I(_1866_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6322__C (.I(_1866_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6286__C (.I(_1866_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5201__C (.I(_1866_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5204__B (.I(_1869_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6961__I1 (.I(_1870_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6490__I3 (.I(_1870_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5954__A2 (.I(_1870_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5206__A1 (.I(_1870_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5463__S (.I(_1873_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5325__S (.I(_1873_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5324__S (.I(_1873_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5209__S (.I(_1873_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5633__I (.I(_1875_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5388__A1 (.I(_1875_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5292__A1 (.I(_1875_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5211__S (.I(_1875_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6261__A2 (.I(_1876_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5218__I1 (.I(_1876_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5366__S (.I(_1877_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5365__S (.I(_1877_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5327__S (.I(_1877_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5213__S (.I(_1877_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6264__A2 (.I(_1878_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5218__I2 (.I(_1878_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5499__A1 (.I(_1879_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5484__A1 (.I(_1879_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5362__S (.I(_1879_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5215__S (.I(_1879_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6262__A2 (.I(_1880_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5218__I3 (.I(_1880_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6381__S (.I(_1881_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5367__S0 (.I(_1881_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5328__S0 (.I(_1881_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5218__S0 (.I(_1881_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5335__S1 (.I(_1882_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5328__S1 (.I(_1882_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5231__S1 (.I(_1882_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5218__S1 (.I(_1882_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5220__A2 (.I(_1883_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6461__A2 (.I(_1886_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5361__A2 (.I(_1886_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5330__A2 (.I(_1886_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5222__A2 (.I(_1886_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6267__I0 (.I(_1889_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5231__I0 (.I(_1889_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5478__S (.I(_1890_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5371__S (.I(_1890_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5268__I (.I(_1890_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5226__S (.I(_1890_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6267__I1 (.I(_1891_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5231__I1 (.I(_1891_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5372__S (.I(_1892_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5333__S (.I(_1892_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5332__S (.I(_1892_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5228__S (.I(_1892_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6270__I1 (.I(_1893_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5231__I2 (.I(_1893_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5906__I (.I(_1894_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5373__S (.I(_1894_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5334__S (.I(_1894_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5230__S (.I(_1894_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6270__I0 (.I(_1895_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5231__I3 (.I(_1895_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5232__A2 (.I(_1896_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5235__B2 (.I(_1897_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6343__C (.I(_1898_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6214__A1 (.I(_1898_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6174__A1 (.I(_1898_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5234__A1 (.I(_1898_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7539__I1 (.I(_1901_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6499__I3 (.I(_1901_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5925__I1 (.I(_1901_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5237__A1 (.I(_1901_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5804__I (.I(_1903_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5379__S (.I(_1903_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5351__A1 (.I(_1903_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5239__S (.I(_1903_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6274__A2 (.I(_1904_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5246__I0 (.I(_1904_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5380__S (.I(_1906_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5341__S (.I(_1906_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5255__A1 (.I(_1906_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5242__S (.I(_1906_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6279__A2 (.I(_1907_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5246__I2 (.I(_1907_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5474__S (.I(_1908_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5381__S (.I(_1908_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5342__S (.I(_1908_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5244__S (.I(_1908_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6197__A1 (.I(_1910_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6155__A1 (.I(_1910_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5343__S0 (.I(_1910_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5246__S0 (.I(_1910_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5247__A2 (.I(_1911_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6380__S0 (.I(_1915_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5558__B2 (.I(_1915_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5529__I (.I(_1915_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5251__S1 (.I(_1915_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5252__A2 (.I(_1916_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5260__A1 (.I(_1917_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5899__S0 (.I(_1918_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5814__S (.I(_1918_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5389__A1 (.I(_1918_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5256__A1 (.I(_1918_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7624__A1 (.I(_1919_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5922__A2 (.I(_1919_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5256__A2 (.I(_1919_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6284__I0 (.I(_1921_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5259__A2 (.I(_1921_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6284__I1 (.I(_1922_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5258__A2 (.I(_1922_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5261__B (.I(_1925_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5265__I (.I(_1929_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6241__A1 (.I(_1931_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6237__A1 (.I(_1931_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6224__A1 (.I(_1931_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5275__A1 (.I(_1931_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6341__S1 (.I(_1932_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5875__S (.I(_1932_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5723__A1 (.I(_1932_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5272__A1 (.I(_1932_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6428__A1 (.I(_1933_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5977__A1 (.I(_1933_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5352__A1 (.I(_1933_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5271__A1 (.I(_1933_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5983__A2 (.I(_1934_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5271__A2 (.I(_1934_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6320__A2 (.I(_1936_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5275__A2 (.I(_1936_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6319__A2 (.I(_1937_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5274__A2 (.I(_1937_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5284__A2 (.I(_1939_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5620__A1 (.I(_1940_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5613__A1 (.I(_1940_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5606__A1 (.I(_1940_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5277__I (.I(_1940_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6366__A1 (.I(_1941_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6338__A1 (.I(_1941_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6274__A1 (.I(_1941_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5280__A1 (.I(_1941_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5520__I (.I(_1942_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5308__A1 (.I(_1942_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5281__S (.I(_1942_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5279__S (.I(_1942_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5284__A3 (.I(_1947_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6312__A2 (.I(_1950_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5295__I0 (.I(_1950_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5765__S (.I(_1951_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5472__A1 (.I(_1951_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5449__A1 (.I(_1951_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5288__S (.I(_1951_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6313__A2 (.I(_1952_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5295__I1 (.I(_1952_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5609__A1 (.I(_1953_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5602__A1 (.I(_1953_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5593__A1 (.I(_1953_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5290__I (.I(_1953_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5863__S (.I(_1954_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5827__S (.I(_1954_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5761__A1 (.I(_1954_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5293__A1 (.I(_1954_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6844__A1 (.I(_1955_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6523__A2 (.I(_1955_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5293__A2 (.I(_1955_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6316__A2 (.I(_1957_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5295__I2 (.I(_1957_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6315__A2 (.I(_1958_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5295__I3 (.I(_1958_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5296__A2 (.I(_1959_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6432__A1 (.I(_1965_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6187__B (.I(_1965_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6084__C (.I(_1965_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5302__I (.I(_1965_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6566__A1 (.I(_1966_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6549__A1 (.I(_1966_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6510__A1 (.I(_1966_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5321__A1 (.I(_1966_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6137__B2 (.I(_1968_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5315__S (.I(_1968_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5310__S (.I(_1968_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5305__S (.I(_1968_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6304__A2 (.I(_1970_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5311__I1 (.I(_1970_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7053__A1 (.I(_1971_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6514__A2 (.I(_1971_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5309__A2 (.I(_1971_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6306__A2 (.I(_1973_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5311__I2 (.I(_1973_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6305__A2 (.I(_1974_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5311__I3 (.I(_1974_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5312__A2 (.I(_1975_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6309__I0 (.I(_1978_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5318__I0 (.I(_1978_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6309__I1 (.I(_1979_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5318__I1 (.I(_1979_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6347__A2 (.I(_1988_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5328__I1 (.I(_1988_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6345__A2 (.I(_1989_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5328__I2 (.I(_1989_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6344__A2 (.I(_1990_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5328__I3 (.I(_1990_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5329__A2 (.I(_1991_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5337__A2 (.I(_1992_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6351__I0 (.I(_1994_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5335__I0 (.I(_1994_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6351__I1 (.I(_1995_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5335__I1 (.I(_1995_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6350__I1 (.I(_1996_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5335__I2 (.I(_1996_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6350__I0 (.I(_1997_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5335__I3 (.I(_1997_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5336__A2 (.I(_1998_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5337__B2 (.I(_1999_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6338__A2 (.I(_2002_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5343__I0 (.I(_2002_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6337__A2 (.I(_2003_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5343__I1 (.I(_2003_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5344__A2 (.I(_2006_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6137__A1 (.I(_2009_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5541__B2 (.I(_2009_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5385__S1 (.I(_2009_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5347__S1 (.I(_2009_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5348__A2 (.I(_2010_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6347__A1 (.I(_2012_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6088__A1 (.I(_2012_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5392__A1 (.I(_2012_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5355__A1 (.I(_2012_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7629__A1 (.I(_2013_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5996__A2 (.I(_2013_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5352__A2 (.I(_2013_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6342__I0 (.I(_2015_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5355__A2 (.I(_2015_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6342__I1 (.I(_2016_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5354__A2 (.I(_2016_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5357__B (.I(_2019_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5360__I (.I(_2022_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6365__A2 (.I(_2024_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5367__I0 (.I(_2024_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5862__S0 (.I(_2025_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5826__S0 (.I(_2025_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5712__I (.I(_2025_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5364__S (.I(_2025_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6367__A2 (.I(_2028_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5367__I3 (.I(_2028_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5368__A2 (.I(_2029_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6370__I0 (.I(_2032_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5374__I0 (.I(_2032_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6371__I1 (.I(_2035_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5374__I3 (.I(_2035_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6374__A2 (.I(_2040_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5383__I0 (.I(_2040_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6373__A2 (.I(_2041_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5383__I1 (.I(_2041_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6351__S (.I(_2044_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6321__S (.I(_2044_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6284__S (.I(_2044_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5383__S0 (.I(_2044_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5384__A2 (.I(_2045_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5386__A2 (.I(_2047_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6381__I0 (.I(_2051_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5392__A2 (.I(_2051_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6381__I1 (.I(_2052_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5391__A2 (.I(_2052_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5394__B (.I(_2055_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5397__I (.I(_2058_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6291__I (.I(_2059_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5500__I (.I(_2059_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5489__I (.I(_2059_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5399__I (.I(_2059_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6532__A1 (.I(_2061_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6017__A1 (.I(_2061_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5580__A1 (.I(_2061_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5401__I (.I(_2061_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6058__A1 (.I(_2062_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6005__A1 (.I(_2062_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5952__A1 (.I(_2062_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5402__I (.I(_2062_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6458__A1 (.I(_2063_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5641__A1 (.I(_2063_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5435__A1 (.I(_2063_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5409__A1 (.I(_2063_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5725__A1 (.I(_2068_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5668__A1 (.I(_2068_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5654__A1 (.I(_2068_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5408__I (.I(_2068_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5682__I (.I(_2069_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5460__A1 (.I(_2069_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5436__I (.I(_2069_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5411__I (.I(_2069_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6245__B2 (.I(_2070_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6184__A1 (.I(_2070_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5565__A1 (.I(_2070_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5412__I (.I(_2070_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6537__A1 (.I(_2071_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6436__A1 (.I(_2071_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5710__A1 (.I(_2071_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5413__I (.I(_2071_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6485__A1 (.I(_2072_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5487__A1 (.I(_2072_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5440__A1 (.I(_2072_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5419__A1 (.I(_2072_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6464__B (.I(_2073_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6444__C (.I(_2073_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6182__A1 (.I(_2073_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5415__I (.I(_2073_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5669__A1 (.I(_2074_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5476__A1 (.I(_2074_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5440__A2 (.I(_2074_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5419__A2 (.I(_2074_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5954__B (.I(_2075_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5630__I (.I(_2075_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5486__A2 (.I(_2075_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5417__I (.I(_2075_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5675__A1 (.I(_2076_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5440__A3 (.I(_2076_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5433__A3 (.I(_2076_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5418__I (.I(_2076_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5441__A2 (.I(_2077_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5434__A2 (.I(_2077_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5423__A2 (.I(_2077_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5419__A3 (.I(_2077_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6372__C (.I(_2078_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6311__C (.I(_2078_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5445__A1 (.I(_2078_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5421__I (.I(_2078_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6528__C (.I(_2079_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6251__A1 (.I(_2079_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5990__A1 (.I(_2079_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5422__I (.I(_2079_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5912__A1 (.I(_2080_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5441__A1 (.I(_2080_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5434__A1 (.I(_2080_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5423__A1 (.I(_2080_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6084__A1 (.I(_2081_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5526__A1 (.I(_2081_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5456__A1 (.I(_2081_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5425__A1 (.I(_2081_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5715__A1 (.I(_2082_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5706__A1 (.I(_2082_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5695__A1 (.I(_2082_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5427__A2 (.I(_2082_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6133__C (.I(_2084_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5640__A1 (.I(_2084_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5502__B (.I(_2084_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5430__I (.I(_2084_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5872__A1 (.I(_2085_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5840__A1 (.I(_2085_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5503__A1 (.I(_2085_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5433__A1 (.I(_2085_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5618__A2 (.I(_2086_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5611__A2 (.I(_2086_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5539__I (.I(_2086_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5432__I (.I(_2086_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6082__A2 (.I(_2087_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6077__A1 (.I(_2087_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5524__A2 (.I(_2087_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5433__A2 (.I(_2087_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5704__B (.I(_2088_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5648__I (.I(_2088_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5584__B2 (.I(_2088_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5437__I (.I(_2088_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6129__B2 (.I(_2089_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5679__A1 (.I(_2089_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5628__A1 (.I(_2089_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5438__A1 (.I(_2089_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6541__A1 (.I(_2091_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6022__C (.I(_2091_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5655__A1 (.I(_2091_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5446__A1 (.I(_2091_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6441__I (.I(_2092_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6417__I (.I(_2092_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6396__I (.I(_2092_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5444__A1 (.I(_2092_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6230__B2 (.I(_2093_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5588__A3 (.I(_2093_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5518__A2 (.I(_2093_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5445__A2 (.I(_2093_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5690__I (.I(_2096_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5564__I (.I(_2096_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5483__I (.I(_2096_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5448__I (.I(_2096_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6033__A1 (.I(_2097_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5921__A1 (.I(_2097_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5473__A1 (.I(_2097_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5450__A1 (.I(_2097_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5776__A2 (.I(_2099_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5628__A2 (.I(_2099_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5467__A2 (.I(_2099_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6405__I (.I(_2100_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5936__B (.I(_2100_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5810__I (.I(_2100_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5455__A1 (.I(_2100_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5873__I (.I(_2101_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5763__I (.I(_2101_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5453__I (.I(_2101_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6551__B (.I(_2103_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6496__A1 (.I(_2103_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6492__B (.I(_2103_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5455__A2 (.I(_2103_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6009__A1 (.I(_2104_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5989__B2 (.I(_2104_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5503__C (.I(_2104_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5456__A2 (.I(_2104_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5862__S1 (.I(_2106_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5826__S1 (.I(_2106_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5752__A1 (.I(_2106_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5458__I (.I(_2106_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6506__I (.I(_2107_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6247__A1 (.I(_2107_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6217__I (.I(_2107_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5459__I (.I(_2107_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6556__C (.I(_2108_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6495__C (.I(_2108_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6248__A1 (.I(_2108_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5462__A1 (.I(_2108_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6406__A1 (.I(_2110_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5797__A1 (.I(_2110_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5482__A1 (.I(_2110_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5462__A2 (.I(_2110_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5738__A1 (.I(_2112_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5638__A2 (.I(_2112_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5466__A2 (.I(_2112_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6094__B2 (.I(_2116_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5895__I (.I(_2116_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5700__A1 (.I(_2116_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5469__A1 (.I(_2116_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6028__A2 (.I(_2118_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5898__A1 (.I(_2118_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5669__A2 (.I(_2118_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5476__A2 (.I(_2118_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5515__A1 (.I(_2119_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5508__A1 (.I(_2119_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5496__A1 (.I(_2119_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5476__B1 (.I(_2119_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5653__A2 (.I(_2121_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5476__B2 (.I(_2121_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5808__A2 (.I(_2122_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5645__A2 (.I(_2122_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5475__A2 (.I(_2122_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5869__A1 (.I(_2124_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5666__A2 (.I(_2124_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5479__A2 (.I(_2124_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5849__A2 (.I(_2125_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5660__A2 (.I(_2125_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5479__B1 (.I(_2125_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5908__A1 (.I(_2127_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5670__A2 (.I(_2127_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5482__A2 (.I(_2127_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6245__A1 (.I(_2129_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6050__A1 (.I(_2129_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5711__A1 (.I(_2129_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5485__A1 (.I(_2129_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5883__A2 (.I(_2131_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5679__A2 (.I(_2131_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5488__B1 (.I(_2131_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5515__B2 (.I(_2133_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5508__B2 (.I(_2133_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5496__B2 (.I(_2133_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5488__B2 (.I(_2133_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6384__A1 (.I(_2134_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6354__A1 (.I(_2134_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6324__A1 (.I(_2134_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5490__I (.I(_2134_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5677__A1 (.I(_2135_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5663__A1 (.I(_2135_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5505__A1 (.I(_2135_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5492__A1 (.I(_2135_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5945__A2 (.I(_2137_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5689__A2 (.I(_2137_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5496__A2 (.I(_2137_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5584__A1 (.I(_2138_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5514__A1 (.I(_2138_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5507__A1 (.I(_2138_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5495__A1 (.I(_2138_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5924__A2 (.I(_2140_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5694__A2 (.I(_2140_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5496__B1 (.I(_2140_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5988__A2 (.I(_2142_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5705__A2 (.I(_2142_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5503__A2 (.I(_2142_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5965__A2 (.I(_2143_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5700__A2 (.I(_2143_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5502__A1 (.I(_2143_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6296__A1 (.I(_2144_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5928__I (.I(_2144_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5509__I (.I(_2144_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5501__A1 (.I(_2144_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5965__A3 (.I(_2145_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5700__A3 (.I(_2145_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5502__A2 (.I(_2145_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6020__A2 (.I(_2148_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5710__A2 (.I(_2148_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5508__A2 (.I(_2148_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5999__A2 (.I(_2150_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5714__A2 (.I(_2150_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5508__B1 (.I(_2150_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6469__A1 (.I(_2151_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5922__A1 (.I(_2151_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5656__A1 (.I(_2151_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5512__A1 (.I(_2151_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5868__S (.I(_2152_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5836__S (.I(_2152_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5812__A1 (.I(_2152_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5511__A1 (.I(_2152_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6053__A2 (.I(_2154_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5721__A2 (.I(_2154_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5515__A2 (.I(_2154_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6036__A2 (.I(_2156_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5724__A2 (.I(_2156_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5515__B1 (.I(_2156_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6329__B1 (.I(_2157_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6298__B1 (.I(_2157_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6139__B1 (.I(_2157_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5517__I (.I(_2157_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5568__A1 (.I(_2159_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5553__B1 (.I(_2159_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5526__B1 (.I(_2159_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6240__A1 (.I(_2160_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6238__A1 (.I(_2160_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6235__A1 (.I(_2160_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5524__B1 (.I(_2160_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5958__S (.I(_2161_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5879__S (.I(_2161_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5853__A1 (.I(_2161_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5522__A1 (.I(_2161_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6105__B2 (.I(_2162_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5951__I (.I(_2162_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5737__I (.I(_2162_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5522__B2 (.I(_2162_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5524__B2 (.I(_2164_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6084__B1 (.I(_2165_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5526__B2 (.I(_2165_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5725__B2 (.I(_2168_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5662__A1 (.I(_2168_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5647__A1 (.I(_2168_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5534__A2 (.I(_2168_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6231__A1 (.I(_2169_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6131__A1 (.I(_2169_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5553__A1 (.I(_2169_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5532__A1 (.I(_2169_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6540__C (.I(_2170_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5869__C2 (.I(_2170_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5837__C2 (.I(_2170_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5531__A1 (.I(_2170_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6490__S1 (.I(_2171_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6467__A1 (.I(_2171_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6409__A1 (.I(_2171_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5531__B2 (.I(_2171_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6071__A1 (.I(_2172_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5532__A2 (.I(_2172_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5534__A3 (.I(_2174_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5622__B2 (.I(_2177_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5615__B2 (.I(_2177_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5608__B2 (.I(_2177_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5538__I (.I(_2177_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5601__B2 (.I(_2178_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5587__B2 (.I(_2178_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5570__A1 (.I(_2178_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5555__A1 (.I(_2178_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5586__A2 (.I(_2179_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5581__A2 (.I(_2179_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5560__A2 (.I(_2179_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5543__A2 (.I(_2179_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6371__S (.I(_2180_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6193__A1 (.I(_2180_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6151__A1 (.I(_2180_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5542__A1 (.I(_2180_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5543__C (.I(_2182_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6132__A1 (.I(_2183_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5555__A2 (.I(_2183_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6476__A1 (.I(_2184_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6420__A1 (.I(_2184_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5569__A1 (.I(_2184_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5554__A1 (.I(_2184_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6110__A1 (.I(_2185_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6053__A1 (.I(_2185_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6020__A1 (.I(_2185_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5553__A2 (.I(_2185_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6209__A1 (.I(_2186_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6169__A1 (.I(_2186_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6102__A1 (.I(_2186_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5551__A1 (.I(_2186_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5755__A1 (.I(_2187_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5731__A1 (.I(_2187_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5616__B2 (.I(_2187_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5548__I (.I(_2187_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6189__B2 (.I(_2188_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6157__B2 (.I(_2188_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6144__B2 (.I(_2188_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5550__A1 (.I(_2188_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6477__I (.I(_2189_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5938__S (.I(_2189_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5558__A1 (.I(_2189_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5550__B2 (.I(_2189_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5552__C (.I(_2191_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6141__A1 (.I(_2192_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5553__B2 (.I(_2192_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6126__A2 (.I(_2195_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6099__A1 (.I(_2195_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5586__B1 (.I(_2195_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5560__B1 (.I(_2195_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6210__A1 (.I(_2196_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6170__A1 (.I(_2196_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6095__A1 (.I(_2196_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5559__A1 (.I(_2196_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6177__A1 (.I(_2199_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5570__A2 (.I(_2199_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6186__A2 (.I(_2200_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6180__A2 (.I(_2200_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6130__A2 (.I(_2200_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5567__A2 (.I(_2200_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6386__B1 (.I(_2201_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6356__B1 (.I(_2201_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6085__A2 (.I(_2201_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5563__I (.I(_2201_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6247__B (.I(_2202_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6186__B1 (.I(_2202_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6180__B1 (.I(_2202_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5567__B1 (.I(_2202_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6501__I (.I(_2203_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6184__B2 (.I(_2203_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5702__A1 (.I(_2203_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5565__B2 (.I(_2203_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6183__A1 (.I(_2206_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5568__A2 (.I(_2206_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6537__A2 (.I(_2210_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6247__C (.I(_2210_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5767__A1 (.I(_2210_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5573__I (.I(_2210_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6545__B2 (.I(_2211_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6505__B2 (.I(_2211_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5904__A1 (.I(_2211_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5582__A1 (.I(_2211_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6250__A1 (.I(_2212_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6218__A1 (.I(_2212_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6082__B1 (.I(_2212_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5582__A2 (.I(_2212_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6047__A1 (.I(_2214_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5995__A1 (.I(_2214_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5967__I (.I(_2214_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5577__A1 (.I(_2214_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6384__B2 (.I(_2216_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6354__B2 (.I(_2216_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5626__I (.I(_2216_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5579__I (.I(_2216_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6225__A1 (.I(_2217_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5723__B (.I(_2217_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5652__B (.I(_2217_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5580__B (.I(_2217_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6218__A2 (.I(_2219_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5582__A3 (.I(_2219_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6246__A2 (.I(_2221_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5607__A2 (.I(_2221_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5600__A2 (.I(_2221_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5585__A1 (.I(_2221_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6248__A2 (.I(_2224_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5587__B1 (.I(_2224_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5622__A1 (.I(_2225_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5615__A1 (.I(_2225_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5608__A1 (.I(_2225_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5601__A1 (.I(_2225_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6278__I (.I(_2228_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5610__A1 (.I(_2228_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5603__A1 (.I(_2228_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5594__A1 (.I(_2228_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6299__I0 (.I(_2232_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5601__A2 (.I(_2232_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5600__C (.I(_2236_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6299__I1 (.I(_2237_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5601__B1 (.I(_2237_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6330__I0 (.I(_2240_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5608__A2 (.I(_2240_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6330__I1 (.I(_2243_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5608__B1 (.I(_2243_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6360__I0 (.I(_2246_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5615__A2 (.I(_2246_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5614__C (.I(_2248_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6360__I1 (.I(_2249_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5615__B1 (.I(_2249_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5618__C (.I(_2251_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6390__I0 (.I(_2252_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5622__A2 (.I(_2252_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6390__I1 (.I(_2255_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5622__B1 (.I(_2255_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6402__A1 (.I(_2256_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5941__A1 (.I(_2256_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5697__A1 (.I(_2256_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5624__A1 (.I(_2256_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6451__A1 (.I(_2258_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6413__S (.I(_2258_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5925__S (.I(_2258_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5627__A1 (.I(_2258_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5699__B (.I(_2259_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5678__B (.I(_2259_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5665__B (.I(_2259_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5627__B (.I(_2259_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6398__A2 (.I(_2261_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5629__A2 (.I(_2261_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6053__C (.I(_2263_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6020__C (.I(_2263_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5966__C (.I(_2263_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5640__A2 (.I(_2263_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6481__A1 (.I(_2264_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5962__A1 (.I(_2264_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5642__A1 (.I(_2264_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5632__A1 (.I(_2264_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5953__A1 (.I(_2266_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5950__A1 (.I(_2266_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5885__A1 (.I(_2266_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5636__A1 (.I(_2266_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6327__B2 (.I(_2267_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6296__B2 (.I(_2267_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5687__I (.I(_2267_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5635__I (.I(_2267_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5673__C (.I(_2268_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5658__B (.I(_2268_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5644__B (.I(_2268_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5636__B (.I(_2268_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6499__S0 (.I(_2270_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5670__A1 (.I(_2270_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5645__A1 (.I(_2270_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5638__A1 (.I(_2270_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6418__A2 (.I(_2272_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5640__A3 (.I(_2272_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6470__A1 (.I(_2275_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6008__S (.I(_2275_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5893__A1 (.I(_2275_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5644__A1 (.I(_2275_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6424__A2 (.I(_2278_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5647__A2 (.I(_2278_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5724__A1 (.I(_2280_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5720__B (.I(_2280_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5694__A1 (.I(_2280_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5653__A1 (.I(_2280_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5856__A1 (.I(_2281_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5817__A1 (.I(_2281_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5722__A1 (.I(_2281_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5650__A1 (.I(_2281_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5960__S (.I(_2283_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5946__I (.I(_2283_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5818__A1 (.I(_2283_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5652__A1 (.I(_2283_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6443__A2 (.I(_2285_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5654__A2 (.I(_2285_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6057__A1 (.I(_2288_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6039__A1 (.I(_2288_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5673__A1 (.I(_2288_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5658__A1 (.I(_2288_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6490__S0 (.I(_2290_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5766__B2 (.I(_2290_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5666__A1 (.I(_2290_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5660__A1 (.I(_2290_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6447__A2 (.I(_2292_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5662__A2 (.I(_2292_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6079__I (.I(_2295_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6059__S (.I(_2295_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5678__A1 (.I(_2295_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5665__A1 (.I(_2295_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6463__A2 (.I(_2298_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5668__A2 (.I(_2298_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6426__A1 (.I(_2301_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5979__A1 (.I(_2301_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5935__S (.I(_2301_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5672__A1 (.I(_2301_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6474__A2 (.I(_2304_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5675__A2 (.I(_2304_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5715__B2 (.I(_2306_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5706__B2 (.I(_2306_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5695__B2 (.I(_2306_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5680__A1 (.I(_2306_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6486__A2 (.I(_2309_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5680__A2 (.I(_2309_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6178__B2 (.I(_2311_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5713__B (.I(_2311_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5693__B (.I(_2311_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5683__I (.I(_2311_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6557__A1 (.I(_2312_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6437__A1 (.I(_2312_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5721__A1 (.I(_2312_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5689__A1 (.I(_2312_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5996__A1 (.I(_2313_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5775__A1 (.I(_2313_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5708__A1 (.I(_2313_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5685__A1 (.I(_2313_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6523__A1 (.I(_2315_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6478__A1 (.I(_2315_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5709__A1 (.I(_2315_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5688__A1 (.I(_2315_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6498__A2 (.I(_2318_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5695__A2 (.I(_2318_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6225__B2 (.I(_2319_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6178__A1 (.I(_2319_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5884__I (.I(_2319_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5691__A1 (.I(_2319_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6522__A1 (.I(_2321_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5902__S (.I(_2321_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5813__A1 (.I(_2321_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5693__A1 (.I(_2321_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6507__A2 (.I(_2323_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5695__B1 (.I(_2323_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6094__A1 (.I(_2326_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6037__S (.I(_2326_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5940__A1 (.I(_2326_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5699__A1 (.I(_2326_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6517__A2 (.I(_2329_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5706__A2 (.I(_2329_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6032__S (.I(_2331_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5997__S (.I(_2331_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5905__S (.I(_2331_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5704__A1 (.I(_2331_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6526__A2 (.I(_2333_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5706__B1 (.I(_2333_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6538__A2 (.I(_2337_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5715__A2 (.I(_2337_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6038__S (.I(_2339_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5926__S (.I(_2339_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5880__S (.I(_2339_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5713__A1 (.I(_2339_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6546__A2 (.I(_2341_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5715__B1 (.I(_2341_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6553__A1 (.I(_2343_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6434__A1 (.I(_2343_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5980__A1 (.I(_2343_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5718__A1 (.I(_2343_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6493__A1 (.I(_2345_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6452__A1 (.I(_2345_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6021__A1 (.I(_2345_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5720__A1 (.I(_2345_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6558__A2 (.I(_2347_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5725__A2 (.I(_2347_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6559__A2 (.I(_2350_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5725__B1 (.I(_2350_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6558__A1 (.I(_2353_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6498__A1 (.I(_2353_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6495__A1 (.I(_2353_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5747__A1 (.I(_2353_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6051__B (.I(_2354_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6018__B (.I(_2354_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5830__I (.I(_2354_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5730__I (.I(_2354_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5847__A1 (.I(_2358_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5806__A1 (.I(_2358_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5740__S (.I(_2358_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5734__S (.I(_2358_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6189__A1 (.I(_2360_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6144__A1 (.I(_2360_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6025__S (.I(_2360_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5736__S (.I(_2360_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6418__C1 (.I(_2361_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5738__C1 (.I(_2361_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5746__A2 (.I(_2364_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6418__B1 (.I(_2365_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5746__B1 (.I(_2365_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6126__A1 (.I(_2366_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5936__A1 (.I(_2366_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5833__I (.I(_2366_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5745__A1 (.I(_2366_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6415__C2 (.I(_2368_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5744__A2 (.I(_2368_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5790__A2 (.I(_2372_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6121__A1 (.I(_2373_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6118__A1 (.I(_2373_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5749__I (.I(_2373_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6253__I (.I(_2374_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6216__C (.I(_2374_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6176__C (.I(_2374_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5790__A3 (.I(_2374_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6068__A2 (.I(_2375_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5751__I (.I(_2375_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6411__I (.I(_2376_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5881__I (.I(_2376_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5766__C (.I(_2376_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5752__A2 (.I(_2376_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6044__A1 (.I(_2379_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6011__A1 (.I(_2379_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5934__A1 (.I(_2379_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5787__A1 (.I(_2379_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6553__B (.I(_2381_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6427__B (.I(_2381_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5976__I (.I(_2381_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5757__I (.I(_2381_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6457__A2 (.I(_2382_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6450__B (.I(_2382_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6410__B (.I(_2382_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5768__A1 (.I(_2382_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6380__S1 (.I(_2383_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6283__S1 (.I(_2383_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5857__A1 (.I(_2383_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5759__S (.I(_2383_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6404__B1 (.I(_2384_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5768__A2 (.I(_2384_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6562__A1 (.I(_2385_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6408__I (.I(_2385_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5978__A1 (.I(_2385_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5762__A1 (.I(_2385_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6406__A2 (.I(_2387_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5767__A2 (.I(_2387_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6430__B2 (.I(_2388_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6423__I (.I(_2388_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6023__I (.I(_2388_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5766__A1 (.I(_2388_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6404__A2 (.I(_2389_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5766__A2 (.I(_2389_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5766__B1 (.I(_2390_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5787__A2 (.I(_2393_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6531__B (.I(_2394_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5988__A1 (.I(_2394_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5914__I (.I(_2394_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5776__A1 (.I(_2394_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5877__I (.I(_2395_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5805__I (.I(_2395_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5771__I (.I(_2395_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5988__B1 (.I(_2397_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5981__B2 (.I(_2397_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5963__A1 (.I(_2397_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5776__B1 (.I(_2397_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5983__A1 (.I(_2398_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5855__S (.I(_2398_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5834__S (.I(_2398_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5774__A1 (.I(_2398_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5776__B2 (.I(_2400_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6064__A2 (.I(_2402_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5937__I (.I(_2402_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5918__I (.I(_2402_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5778__I (.I(_2402_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5987__B2 (.I(_2403_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5849__B2 (.I(_2403_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5808__B2 (.I(_2403_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5780__A1 (.I(_2403_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6398__C1 (.I(_2404_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5780__A2 (.I(_2404_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6523__B (.I(_2406_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6514__B (.I(_2406_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5987__A1 (.I(_2406_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5783__A1 (.I(_2406_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6398__B2 (.I(_2407_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5783__A2 (.I(_2407_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6061__A1 (.I(_2410_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5974__A1 (.I(_2410_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5955__A1 (.I(_2410_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5786__B (.I(_2410_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5790__B1 (.I(_2412_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6063__B2 (.I(_2414_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5991__A1 (.I(_2414_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5957__B2 (.I(_2414_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5790__B2 (.I(_2414_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6027__A1 (.I(_2416_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5897__A1 (.I(_2416_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5861__A1 (.I(_2416_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5822__A1 (.I(_2416_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6552__A1 (.I(_2417_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6435__A1 (.I(_2417_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5843__A1 (.I(_2417_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5796__A1 (.I(_2417_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6401__A1 (.I(_2418_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6012__S (.I(_2418_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5842__A1 (.I(_2418_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5795__A1 (.I(_2418_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6424__B2 (.I(_2420_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5797__A2 (.I(_2420_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6471__A1 (.I(_2422_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6403__A1 (.I(_2422_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5815__I (.I(_2422_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5799__I (.I(_2422_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6042__A1 (.I(_2423_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5932__A1 (.I(_2423_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5883__A1 (.I(_2423_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5808__A1 (.I(_2423_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6530__A1 (.I(_2424_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5984__A1 (.I(_2424_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5846__A1 (.I(_2424_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5803__A1 (.I(_2424_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6199__A1 (.I(_2425_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6157__A1 (.I(_2425_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5845__A1 (.I(_2425_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5802__A1 (.I(_2425_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6424__C1 (.I(_2427_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5808__B1 (.I(_2427_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6030__A1 (.I(_2428_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5916__A1 (.I(_2428_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5848__A1 (.I(_2428_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5807__A1 (.I(_2428_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6422__I (.I(_2429_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6397__I (.I(_2429_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5848__B (.I(_2429_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5807__B (.I(_2429_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5808__C (.I(_2431_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6516__C (.I(_2434_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6043__A1 (.I(_2434_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5933__A1 (.I(_2434_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5821__A1 (.I(_2434_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6035__B2 (.I(_2435_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5923__B2 (.I(_2435_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5859__A1 (.I(_2435_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5820__A1 (.I(_2435_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6430__A2 (.I(_2437_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5820__A2 (.I(_2437_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6493__B (.I(_2440_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5915__I (.I(_2440_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5858__A1 (.I(_2440_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5819__A1 (.I(_2440_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5820__C (.I(_2443_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5821__A2 (.I(_2444_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6538__A1 (.I(_2447_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6424__A1 (.I(_2447_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5866__A1 (.I(_2447_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5832__A1 (.I(_2447_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6341__S0 (.I(_2448_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6283__S0 (.I(_2448_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6199__B2 (.I(_2448_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5825__I (.I(_2448_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6221__S1 (.I(_2449_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5936__C (.I(_2449_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5865__A1 (.I(_2449_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5831__A1 (.I(_2449_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5831__A2 (.I(_2450_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6440__A2 (.I(_2451_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5831__B1 (.I(_2451_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5867__S (.I(_2452_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5864__S (.I(_2452_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5835__S (.I(_2452_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5829__S (.I(_2452_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6443__B2 (.I(_2453_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5831__C1 (.I(_2453_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5837__A1 (.I(_2458_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6437__A2 (.I(_2459_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5837__B2 (.I(_2459_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6443__C1 (.I(_2460_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5837__C1 (.I(_2460_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5840__B (.I(_2463_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6042__B2 (.I(_2464_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5998__A1 (.I(_2464_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5932__B2 (.I(_2464_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5844__A1 (.I(_2464_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6447__B2 (.I(_2466_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5844__A2 (.I(_2466_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6447__C1 (.I(_2469_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5849__B1 (.I(_2469_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5849__C (.I(_2471_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6544__B (.I(_2474_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6536__A1 (.I(_2474_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6504__B (.I(_2474_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5860__A1 (.I(_2474_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6514__A1 (.I(_2475_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6482__A1 (.I(_2475_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5961__A1 (.I(_2475_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5854__A1 (.I(_2475_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6454__C2 (.I(_2477_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5859__A2 (.I(_2477_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6454__A2 (.I(_2478_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5859__B1 (.I(_2478_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5859__C (.I(_2481_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5865__A2 (.I(_2485_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6461__B2 (.I(_2486_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5865__B1 (.I(_2486_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6463__B2 (.I(_2487_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5865__C1 (.I(_2487_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6460__A2 (.I(_2490_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5869__B2 (.I(_2490_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5872__B (.I(_2494_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6559__C2 (.I(_2496_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6517__C2 (.I(_2496_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6443__C2 (.I(_2496_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5876__A1 (.I(_2496_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6486__B2 (.I(_2497_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5876__A2 (.I(_2497_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6453__I (.I(_2499_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6442__I (.I(_2499_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6400__I (.I(_2499_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5878__I (.I(_2499_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6546__B1 (.I(_2500_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6524__A1 (.I(_2500_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6507__B1 (.I(_2500_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5882__A1 (.I(_2500_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5882__A2 (.I(_2501_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6486__C1 (.I(_2502_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5882__B1 (.I(_2502_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6564__A1 (.I(_2503_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6454__A1 (.I(_2503_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6404__B2 (.I(_2503_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5882__B2 (.I(_2503_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5898__A2 (.I(_2505_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6031__A1 (.I(_2506_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5954__A1 (.I(_2506_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5917__A1 (.I(_2506_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5887__A1 (.I(_2506_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6557__A2 (.I(_2508_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6526__A1 (.I(_2508_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6218__B (.I(_2508_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5887__C (.I(_2508_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6485__A2 (.I(_2509_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5897__A2 (.I(_2509_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6474__C2 (.I(_2510_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6398__C2 (.I(_2510_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5973__A1 (.I(_2510_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5896__A1 (.I(_2510_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6551__A1 (.I(_2511_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6492__A1 (.I(_2511_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5894__A1 (.I(_2511_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5892__A1 (.I(_2511_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6438__S (.I(_2512_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6014__A1 (.I(_2512_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5930__A1 (.I(_2512_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5891__A1 (.I(_2512_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6484__A2 (.I(_2514_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5896__A2 (.I(_2514_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5896__B1 (.I(_2516_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6080__B2 (.I(_2517_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6066__A1 (.I(_2517_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5903__A1 (.I(_2517_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5896__B2 (.I(_2517_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5912__A2 (.I(_2520_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5903__A2 (.I(_2521_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6539__A1 (.I(_2522_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6533__A1 (.I(_2522_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5982__S (.I(_2522_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5901__S (.I(_2522_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6474__B2 (.I(_2523_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5903__B1 (.I(_2523_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6472__B1 (.I(_2524_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5903__C1 (.I(_2524_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6472__A2 (.I(_2527_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5908__B2 (.I(_2527_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6513__A1 (.I(_2528_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6024__S (.I(_2528_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5972__S (.I(_2528_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5907__S (.I(_2528_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6474__C1 (.I(_2529_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5908__C1 (.I(_2529_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6062__A1 (.I(_2531_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5975__A1 (.I(_2531_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5956__A1 (.I(_2531_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5910__B (.I(_2531_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5912__B (.I(_2533_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6529__A1 (.I(_2534_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6252__A1 (.I(_2534_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6063__A1 (.I(_2534_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5957__A1 (.I(_2534_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6498__B1 (.I(_2536_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6461__B1 (.I(_2536_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6036__B1 (.I(_2536_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5924__B1 (.I(_2536_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5924__B2 (.I(_2538_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6052__A1 (.I(_2539_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6035__A1 (.I(_2539_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5998__B2 (.I(_2539_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5923__A1 (.I(_2539_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6112__A1 (.I(_2540_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6045__S (.I(_2540_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5971__S (.I(_2540_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5920__S (.I(_2540_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6507__C1 (.I(_2541_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5923__A2 (.I(_2541_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6507__B2 (.I(_2543_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5923__B1 (.I(_2543_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6505__A2 (.I(_2547_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5932__B1 (.I(_2547_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6554__A1 (.I(_2548_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6041__A1 (.I(_2548_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6015__A1 (.I(_2548_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5931__A1 (.I(_2548_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6040__A1 (.I(_2549_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6034__A1 (.I(_2549_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6013__A1 (.I(_2549_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5929__A1 (.I(_2549_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5932__C (.I(_2552_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5933__A2 (.I(_2553_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5957__A2 (.I(_2555_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6498__B2 (.I(_2556_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5936__A2 (.I(_2556_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6525__A1 (.I(_2558_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6019__A1 (.I(_2558_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5964__A1 (.I(_2558_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5943__A1 (.I(_2558_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6496__A2 (.I(_2559_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5943__A2 (.I(_2559_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6430__A1 (.I(_2560_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6048__A1 (.I(_2560_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5992__I (.I(_2560_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5942__A1 (.I(_2560_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5943__B (.I(_2563_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6060__A1 (.I(_2565_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6026__B2 (.I(_2565_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5973__B2 (.I(_2565_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5945__C (.I(_2565_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6521__A1 (.I(_2567_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6219__A1 (.I(_2567_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6066__B2 (.I(_2567_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5949__A1 (.I(_2567_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6546__C2 (.I(_2568_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6507__C2 (.I(_2568_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6454__B2 (.I(_2568_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5949__B (.I(_2568_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5955__A2 (.I(_2570_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6219__A2 (.I(_2572_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6058__C (.I(_2572_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5970__C (.I(_2572_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5952__C (.I(_2572_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5955__A3 (.I(_2573_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5956__A3 (.I(_2576_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6517__B2 (.I(_2578_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5959__A2 (.I(_2578_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5966__A1 (.I(_2579_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6517__C1 (.I(_2580_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5964__A2 (.I(_2580_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5964__B (.I(_2583_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6511__A1 (.I(_2587_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6022__A1 (.I(_2587_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5994__A1 (.I(_2587_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5970__A1 (.I(_2587_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6221__S0 (.I(_2588_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6004__A1 (.I(_2588_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5993__A1 (.I(_2588_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5969__A1 (.I(_2588_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5974__A2 (.I(_2590_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6515__A2 (.I(_2591_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5973__A2 (.I(_2591_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5975__A3 (.I(_2594_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6561__A2 (.I(_2596_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6521__B (.I(_2596_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6512__B (.I(_2596_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5981__A1 (.I(_2596_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5978__B (.I(_2597_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6525__A2 (.I(_2598_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5981__A2 (.I(_2598_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5981__B1 (.I(_2600_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6524__A2 (.I(_2602_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5989__B1 (.I(_2602_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5988__B2 (.I(_2604_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6526__B2 (.I(_2605_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5987__A2 (.I(_2605_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6526__C1 (.I(_2606_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5987__B1 (.I(_2606_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5988__C (.I(_2607_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5990__A2 (.I(_2609_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6545__A1 (.I(_2611_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6505__A1 (.I(_2611_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6006__B2 (.I(_2611_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5999__B1 (.I(_2611_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5999__B2 (.I(_2613_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6546__B2 (.I(_2615_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5998__A2 (.I(_2615_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6546__C1 (.I(_2616_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5998__B1 (.I(_2616_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6011__A2 (.I(_2618_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6540__A1 (.I(_2619_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6459__A1 (.I(_2619_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6129__A1 (.I(_2619_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6003__A1 (.I(_2619_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6429__A1 (.I(_2620_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6105__A1 (.I(_2620_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6046__A1 (.I(_2620_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6002__A1 (.I(_2620_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6003__B (.I(_2621_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6541__A2 (.I(_2622_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6006__A2 (.I(_2622_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6006__B1 (.I(_2624_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6011__B1 (.I(_2625_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6528__A1 (.I(_2626_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6433__A1 (.I(_2626_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6419__A1 (.I(_2626_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6011__B2 (.I(_2626_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6545__A2 (.I(_2627_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6009__A2 (.I(_2627_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6538__B1 (.I(_2631_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6019__A2 (.I(_2631_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6019__B (.I(_2634_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6537__A3 (.I(_2636_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6018__A2 (.I(_2636_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6020__B (.I(_2638_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6027__A2 (.I(_2641_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6558__B2 (.I(_2642_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6538__B2 (.I(_2642_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6457__B1 (.I(_2642_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6026__A1 (.I(_2642_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6535__A2 (.I(_2643_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6026__A2 (.I(_2643_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6028__A4 (.I(_2646_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6036__B2 (.I(_2649_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6559__C1 (.I(_2650_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6035__A2 (.I(_2650_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6559__B2 (.I(_2652_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6035__B1 (.I(_2652_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6564__A2 (.I(_2655_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6042__A2 (.I(_2655_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6564__B1 (.I(_2656_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6042__B1 (.I(_2656_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6042__C (.I(_2659_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6043__A2 (.I(_2660_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6063__A2 (.I(_2662_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6558__B1 (.I(_2663_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6052__A2 (.I(_2663_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6052__B (.I(_2666_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6557__A3 (.I(_2668_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6051__A2 (.I(_2668_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6486__C2 (.I(_2672_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6440__B2 (.I(_2672_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6418__C2 (.I(_2672_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6056__A1 (.I(_2672_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6554__A2 (.I(_2673_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6056__A2 (.I(_2673_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6061__A3 (.I(_2676_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6062__A3 (.I(_2679_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6202__A1 (.I(_2681_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6161__A1 (.I(_2681_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6072__I (.I(_2681_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6065__I (.I(_2681_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6183__A2 (.I(_2682_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6177__A2 (.I(_2682_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6133__A1 (.I(_2682_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6067__A1 (.I(_2682_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6223__A2 (.I(_2685_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6134__I (.I(_2685_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6074__I (.I(_2685_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6069__I (.I(_2685_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6273__I (.I(_2686_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6256__I (.I(_2686_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6213__C (.I(_2686_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6070__I (.I(_2686_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6187__A1 (.I(_2687_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6181__A1 (.I(_2687_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6118__A2 (.I(_2687_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6071__A2 (.I(_2687_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6141__A2 (.I(_2689_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6132__A2 (.I(_2689_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6100__A2 (.I(_2689_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6073__A2 (.I(_2689_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6208__C (.I(_2692_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6168__C (.I(_2692_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6109__A1 (.I(_2692_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6076__A2 (.I(_2692_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6512__A1 (.I(_2696_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6450__A1 (.I(_2696_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6125__A1 (.I(_2696_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6080__A1 (.I(_2696_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6563__C (.I(_2698_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6537__B (.I(_2698_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6395__I (.I(_2698_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6082__C (.I(_2698_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6087__A1 (.I(_2700_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6254__I (.I(_2702_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6227__A2 (.I(_2702_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6086__I (.I(_2702_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6300__A1 (.I(_2703_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6188__B (.I(_2703_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6142__A1 (.I(_2703_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6087__B (.I(_2703_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6260__I (.I(_2706_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6149__I (.I(_2706_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6122__I (.I(_2706_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6090__I (.I(_2706_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6207__A1 (.I(_2708_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6167__A1 (.I(_2708_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6114__C (.I(_2708_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6093__A2 (.I(_2708_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6159__I (.I(_2713_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6147__I (.I(_2713_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6097__I (.I(_2713_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6365__B (.I(_2715_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6264__B (.I(_2715_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6108__C (.I(_2715_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6099__C (.I(_2715_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6317__A1 (.I(_2718_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6280__A1 (.I(_2718_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6235__B (.I(_2718_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6104__A1 (.I(_2718_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6309__S (.I(_2723_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6267__S (.I(_2723_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6234__A1 (.I(_2723_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6107__A1 (.I(_2723_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6110__A3 (.I(_2726_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6550__A1 (.I(_2728_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6491__A1 (.I(_2728_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6427__A1 (.I(_2728_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6113__A1 (.I(_2728_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6378__A1 (.I(_2733_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6241__B (.I(_2733_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6120__C (.I(_2733_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6117__C (.I(_2733_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6125__B1 (.I(_2737_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6242__B (.I(_2738_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6236__B (.I(_2738_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6124__A1 (.I(_2738_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6347__B (.I(_2739_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6210__B (.I(_2739_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6170__B (.I(_2739_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6123__C (.I(_2739_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6125__B2 (.I(_2741_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6243__B (.I(_2743_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6215__C (.I(_2743_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6175__C (.I(_2743_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6127__C (.I(_2743_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6128__B (.I(_2744_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6133__A2 (.I(_2747_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6390__S1 (.I(_2750_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6360__S1 (.I(_2750_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6173__C (.I(_2750_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6140__A1 (.I(_2750_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6359__A2 (.I(_2751_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6329__A2 (.I(_2751_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6298__A2 (.I(_2751_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6139__A2 (.I(_2751_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6358__A1 (.I(_2752_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6328__A1 (.I(_2752_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6297__A1 (.I(_2752_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6138__A1 (.I(_2752_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6140__A2 (.I(_2755_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6330__S1 (.I(_2759_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6299__S1 (.I(_2759_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6195__A1 (.I(_2759_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6153__A1 (.I(_2759_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6345__B (.I(_2763_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6306__B (.I(_2763_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6191__C (.I(_2763_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6148__C (.I(_2763_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6212__B (.I(_2775_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6201__C (.I(_2775_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6172__B (.I(_2775_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6160__C (.I(_2775_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6175__A2 (.I(_2778_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6375__A1 (.I(_2779_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6339__A1 (.I(_2779_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6208__A1 (.I(_2779_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6168__A1 (.I(_2779_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6174__A2 (.I(_2789_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6176__B (.I(_2791_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6181__A2 (.I(_2795_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6187__A2 (.I(_2801_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6215__A2 (.I(_2818_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6214__A2 (.I(_2828_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6216__B (.I(_2830_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6560__A1 (.I(_2831_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6464__A1 (.I(_2831_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6444__B2 (.I(_2831_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6230__A1 (.I(_2831_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6220__A1 (.I(_2832_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6220__A2 (.I(_2833_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6230__B1 (.I(_2835_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6285__I (.I(_2837_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6271__I (.I(_2837_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6224__C (.I(_2837_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6229__A1 (.I(_2838_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6228__C (.I(_2841_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6230__C (.I(_2843_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6336__A1 (.I(_2846_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6276__A1 (.I(_2846_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6239__A1 (.I(_2846_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6233__B (.I(_2846_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6249__B (.I(_2862_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6252__B1 (.I(_2863_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6369__A1 (.I(_2869_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6349__A1 (.I(_2869_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6308__A1 (.I(_2869_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6266__A1 (.I(_2869_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6334__A1 (.I(_2870_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6312__A1 (.I(_2870_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6303__A1 (.I(_2870_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6258__A1 (.I(_2870_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6377__A1 (.I(_2872_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6315__A1 (.I(_2872_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6275__A1 (.I(_2872_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6261__A1 (.I(_2872_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6367__B (.I(_2873_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6313__B (.I(_2873_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6304__B (.I(_2873_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6261__B (.I(_2873_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6365__A1 (.I(_2876_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6346__A1 (.I(_2876_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6306__A1 (.I(_2876_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6264__A1 (.I(_2876_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6282__I (.I(_2881_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6269__I (.I(_2881_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6287__A2 (.I(_2885_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6379__A1 (.I(_2886_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6340__A1 (.I(_2886_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6318__A1 (.I(_2886_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6281__A1 (.I(_2886_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6376__A1 (.I(_2891_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6374__A1 (.I(_2891_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6316__A1 (.I(_2891_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6279__A1 (.I(_2891_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6286__A2 (.I(_2896_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6286__B1 (.I(_2897_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6287__B2 (.I(_2899_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6301__A2 (.I(_2900_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6387__A1 (.I(_2904_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6357__A1 (.I(_2904_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6327__A1 (.I(_2904_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6293__A1 (.I(_2904_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6300__A2 (.I(_2912_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6318__A3 (.I(_2929_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6322__A2 (.I(_2932_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6322__B1 (.I(_2933_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6332__A2 (.I(_2935_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6353__A1 (.I(_2951_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6343__A2 (.I(_2952_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6362__A2 (.I(_2964_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6383__B1 (.I(_2989_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6382__A2 (.I(_2990_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6382__B1 (.I(_2991_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6383__B2 (.I(_2992_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6392__A2 (.I(_2993_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6390__I2 (.I(_2996_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6393__A2 (.I(_3002_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6567__A1 (.I(_3003_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6488__A1 (.I(_3003_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6456__A1 (.I(_3003_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6407__A1 (.I(_3003_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6487__A1 (.I(_3004_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6475__A1 (.I(_3004_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6448__A1 (.I(_3004_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6399__A1 (.I(_3004_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6559__A1 (.I(_3005_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6463__A1 (.I(_3005_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6447__A1 (.I(_3005_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6398__A1 (.I(_3005_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6474__B1 (.I(_3006_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6447__B1 (.I(_3006_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6418__B2 (.I(_3006_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6398__B1 (.I(_3006_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6399__A2 (.I(_3007_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6472__B2 (.I(_3009_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6463__B1 (.I(_3009_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6415__C1 (.I(_3009_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6404__A1 (.I(_3009_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6403__A2 (.I(_3010_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6473__A1 (.I(_3014_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6455__C (.I(_3014_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6416__A1 (.I(_3014_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6406__C (.I(_3014_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6407__A3 (.I(_3015_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6565__A1 (.I(_3017_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6468__A1 (.I(_3017_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6449__A1 (.I(_3017_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6410__A1 (.I(_3017_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6535__B2 (.I(_3020_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6515__B2 (.I(_3020_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6425__A1 (.I(_3020_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6412__I (.I(_3020_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6556__A1 (.I(_3021_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6472__A1 (.I(_3021_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6460__A1 (.I(_3021_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6415__A1 (.I(_3021_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6415__B1 (.I(_3022_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6561__B1 (.I(_3023_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6463__C2 (.I(_3023_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6447__C2 (.I(_3023_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6415__B2 (.I(_3023_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6420__A2 (.I(_3025_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6486__A1 (.I(_3026_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6474__A1 (.I(_3026_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6437__C (.I(_3026_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6418__A1 (.I(_3026_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6419__A2 (.I(_3027_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6486__B1 (.I(_3030_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6484__A1 (.I(_3030_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6440__A1 (.I(_3030_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6424__B1 (.I(_3030_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6480__A1 (.I(_3031_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6468__B (.I(_3031_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6460__B2 (.I(_3031_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6424__C2 (.I(_3031_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6433__A2 (.I(_3032_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6430__B1 (.I(_3037_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6432__A2 (.I(_3039_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6437__B (.I(_3044_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6440__B1 (.I(_3046_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6497__A1 (.I(_3047_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6480__B (.I(_3047_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6460__C (.I(_3047_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6440__C (.I(_3047_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6444__A2 (.I(_3048_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6546__A1 (.I(_3049_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6517__A1 (.I(_3049_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6507__A1 (.I(_3049_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6443__A1 (.I(_3049_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6564__B2 (.I(_3050_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6559__B1 (.I(_3050_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6517__B1 (.I(_3050_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6443__B1 (.I(_3050_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6448__A2 (.I(_3054_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6454__B1 (.I(_3059_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6535__A1 (.I(_3060_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6526__B1 (.I(_3060_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6515__A1 (.I(_3060_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6454__C1 (.I(_3060_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6456__A3 (.I(_3062_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6466__A1 (.I(_3063_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6458__A2 (.I(_3064_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6465__A2 (.I(_3069_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6464__A2 (.I(_3070_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6472__C (.I(_3077_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6476__A2 (.I(_3079_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6475__A2 (.I(_3080_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6542__A1 (.I(_3083_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6500__A1 (.I(_3083_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6499__S1 (.I(_3083_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6479__A1 (.I(_3083_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6480__A2 (.I(_3085_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6484__B (.I(_3089_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6487__A2 (.I(_3092_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6495__A2 (.I(_3095_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6495__B (.I(_3099_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6505__B1 (.I(_3104_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6543__A1 (.I(_3106_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6531__A1 (.I(_3106_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6520__A1 (.I(_3106_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6503__A1 (.I(_3106_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6563__B1 (.I(_3107_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6543__B (.I(_3107_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6526__C2 (.I(_3107_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6503__B (.I(_3107_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6510__B1 (.I(_3110_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6508__A2 (.I(_3112_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6515__C (.I(_3118_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6519__A1 (.I(_3120_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6518__A2 (.I(_3121_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6524__B (.I(_3127_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6528__A2 (.I(_3129_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6527__A2 (.I(_3130_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6535__C (.I(_3137_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6536__A3 (.I(_3138_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6545__C (.I(_3147_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6555__A2 (.I(_3153_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6567__A2 (.I(_3158_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6563__B2 (.I(_3164_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6566__A3 (.I(_3167_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7839__I (.I(_3169_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7822__A2 (.I(_3169_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6572__A2 (.I(_3169_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6569__A2 (.I(_3169_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7829__A1 (.I(_3174_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6576__I (.I(_3174_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6590__A4 (.I(_3179_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6587__A3 (.I(_3179_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6584__A2 (.I(_3179_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6582__A2 (.I(_3179_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6903__I0 (.I(_3228_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6832__I0 (.I(_3228_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6737__I0 (.I(_3228_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6684__I0 (.I(_3228_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7744__A2 (.I(_3232_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7549__A1 (.I(_3232_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7283__A1 (.I(_3232_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6682__A2 (.I(_3232_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7038__I (.I(_3234_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6991__I (.I(_3234_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6732__I (.I(_3234_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6681__I (.I(_3234_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6700__I (.I(_3236_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6683__I (.I(_3236_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6696__S (.I(_3237_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6692__S (.I(_3237_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6688__S (.I(_3237_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6684__S (.I(_3237_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7150__I (.I(_3239_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7017__I (.I(_3239_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6928__I (.I(_3239_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6687__I (.I(_3239_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6905__I0 (.I(_3240_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6834__I0 (.I(_3240_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6739__I0 (.I(_3240_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6688__I0 (.I(_3240_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7153__I (.I(_3242_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7020__I (.I(_3242_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6931__I (.I(_3242_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6691__I (.I(_3242_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6907__I0 (.I(_3243_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6837__I0 (.I(_3243_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6741__I0 (.I(_3243_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6692__I0 (.I(_3243_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7156__I (.I(_3245_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7023__I (.I(_3245_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6934__I (.I(_3245_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6695__I (.I(_3245_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6909__I0 (.I(_3246_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6839__I0 (.I(_3246_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6743__I0 (.I(_3246_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6696__I0 (.I(_3246_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6912__I0 (.I(_3249_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6841__I0 (.I(_3249_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6746__I0 (.I(_3249_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6701__I0 (.I(_3249_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7220__I (.I(_3252_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7119__I (.I(_3252_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6963__I (.I(_3252_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6704__I (.I(_3252_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6941__I0 (.I(_3253_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6914__I0 (.I(_3253_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6748__I0 (.I(_3253_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6705__I0 (.I(_3253_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7165__I (.I(_3255_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7032__I (.I(_3255_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6943__I (.I(_3255_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6708__I (.I(_3255_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6916__I0 (.I(_3256_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6845__I0 (.I(_3256_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6750__I0 (.I(_3256_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6709__I0 (.I(_3256_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7168__I (.I(_3258_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7035__I (.I(_3258_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6946__I (.I(_3258_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6712__I (.I(_3258_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6918__I0 (.I(_3259_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6847__I0 (.I(_3259_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6752__I0 (.I(_3259_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6713__I0 (.I(_3259_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6745__I (.I(_3273_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6736__I (.I(_3273_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6743__S (.I(_3274_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6741__S (.I(_3274_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6739__S (.I(_3274_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6737__S (.I(_3274_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6752__S (.I(_3279_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6750__S (.I(_3279_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6748__S (.I(_3279_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6746__S (.I(_3279_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7569__I (.I(_3292_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7484__I (.I(_3292_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7281__I (.I(_3292_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6771__I (.I(_3292_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7784__I0 (.I(_3293_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7765__I0 (.I(_3293_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7248__I1 (.I(_3293_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6779__I1 (.I(_3293_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7782__A1 (.I(_3294_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7246__A1 (.I(_3294_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7187__A1 (.I(_3294_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6777__A1 (.I(_3294_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7611__A1 (.I(_3296_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7329__A2 (.I(_3296_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7246__A3 (.I(_3296_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6777__A2 (.I(_3296_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7463__I (.I(_3297_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7328__I (.I(_3297_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7282__I (.I(_3297_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6776__I (.I(_3297_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6791__S (.I(_3300_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6787__S (.I(_3300_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6783__S (.I(_3300_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6779__S (.I(_3300_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7786__I0 (.I(_3303_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7767__I0 (.I(_3303_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7250__I1 (.I(_3303_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6783__I1 (.I(_3303_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7533__I (.I(_3305_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7336__I (.I(_3305_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7292__I (.I(_3305_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6786__I (.I(_3305_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7788__I0 (.I(_3306_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7769__I0 (.I(_3306_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7252__I1 (.I(_3306_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6787__I1 (.I(_3306_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7558__I (.I(_3308_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7472__I (.I(_3308_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7196__I (.I(_3308_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6790__I (.I(_3308_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7793__I0 (.I(_3312_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7623__A1 (.I(_3312_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7257__I1 (.I(_3312_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6796__I1 (.I(_3312_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7259__I1 (.I(_3316_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7052__A1 (.I(_3316_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6843__A1 (.I(_3316_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6800__I1 (.I(_3316_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7586__I (.I(_3318_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7501__I (.I(_3318_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7302__I (.I(_3318_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6803__I (.I(_3318_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7797__I0 (.I(_3319_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7628__A1 (.I(_3319_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7261__I1 (.I(_3319_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6804__I1 (.I(_3319_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7589__I (.I(_3321_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7504__I (.I(_3321_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7305__I (.I(_3321_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6807__I (.I(_3321_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7799__I0 (.I(_3322_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7630__A1 (.I(_3322_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7263__I1 (.I(_3322_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6808__I1 (.I(_3322_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7570__A2 (.I(_3335_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7187__A3 (.I(_3335_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7039__A3 (.I(_3335_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6830__A3 (.I(_3335_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6847__S (.I(_3336_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6836__I (.I(_3336_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6831__I (.I(_3336_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6844__A2 (.I(_3337_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6843__A2 (.I(_3337_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6834__S (.I(_3337_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6832__S (.I(_3337_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6845__S (.I(_3340_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6841__S (.I(_3340_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6839__S (.I(_3340_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6837__S (.I(_3340_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7763__A3 (.I(_3371_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7485__A2 (.I(_3371_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6992__A2 (.I(_3371_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6901__A2 (.I(_3371_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6911__I (.I(_3375_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6902__I (.I(_3375_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6909__S (.I(_3376_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6907__S (.I(_3376_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6905__S (.I(_3376_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6903__S (.I(_3376_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6918__S (.I(_3381_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6916__S (.I(_3381_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6914__S (.I(_3381_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6912__S (.I(_3381_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6994__I0 (.I(_3386_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6974__I0 (.I(_3386_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6952__I0 (.I(_3386_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6926__I0 (.I(_3386_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6938__I (.I(_3390_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6925__I (.I(_3390_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6935__S (.I(_3391_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6932__S (.I(_3391_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6929__S (.I(_3391_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6926__S (.I(_3391_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6996__I0 (.I(_3393_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6976__I0 (.I(_3393_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6954__I0 (.I(_3393_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6929__I0 (.I(_3393_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6998__I0 (.I(_3395_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6978__I0 (.I(_3395_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6956__I0 (.I(_3395_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6932__I0 (.I(_3395_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7003__I0 (.I(_3399_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6983__I0 (.I(_3399_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6961__I0 (.I(_3399_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6939__I0 (.I(_3399_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6947__S (.I(_3400_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6944__S (.I(_3400_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6941__S (.I(_3400_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6939__S (.I(_3400_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7007__I0 (.I(_3403_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6987__I0 (.I(_3403_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6966__I0 (.I(_3403_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6944__I0 (.I(_3403_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7009__I0 (.I(_3405_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6989__I0 (.I(_3405_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6968__I0 (.I(_3405_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6947__I0 (.I(_3405_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6960__I (.I(_3408_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6951__I (.I(_3408_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6968__S (.I(_3414_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6966__S (.I(_3414_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6964__S (.I(_3414_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6961__S (.I(_3414_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7030__I0 (.I(_3416_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7005__I0 (.I(_3416_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6985__I0 (.I(_3416_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6964__I0 (.I(_3416_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6982__I (.I(_3422_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6973__I (.I(_3422_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6980__S (.I(_3423_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6978__S (.I(_3423_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6976__S (.I(_3423_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6974__S (.I(_3423_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6989__S (.I(_3428_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6987__S (.I(_3428_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6985__S (.I(_3428_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6983__S (.I(_3428_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7002__I (.I(_3434_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6993__I (.I(_3434_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7000__S (.I(_3435_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6998__S (.I(_3435_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6996__S (.I(_3435_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6994__S (.I(_3435_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7009__S (.I(_3440_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7007__S (.I(_3440_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7005__S (.I(_3440_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7003__S (.I(_3440_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7128__I0 (.I(_3445_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7108__I0 (.I(_3445_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7041__I0 (.I(_3445_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7015__I0 (.I(_3445_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7782__A3 (.I(_3446_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7592__A2 (.I(_3446_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7308__A3 (.I(_3446_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7013__A2 (.I(_3446_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7027__I (.I(_3447_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7014__I (.I(_3447_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7024__S (.I(_3448_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7021__S (.I(_3448_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7018__S (.I(_3448_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7015__S (.I(_3448_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7130__I0 (.I(_3450_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7110__I0 (.I(_3450_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7043__I0 (.I(_3450_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7018__I0 (.I(_3450_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7132__I0 (.I(_3452_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7112__I0 (.I(_3452_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7046__I0 (.I(_3452_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7021__I0 (.I(_3452_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7134__I0 (.I(_3454_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7114__I0 (.I(_3454_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7048__I0 (.I(_3454_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7024__I0 (.I(_3454_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7137__I0 (.I(_3456_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7117__I0 (.I(_3456_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7050__I0 (.I(_3456_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7028__I0 (.I(_3456_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7036__S (.I(_3457_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7033__S (.I(_3457_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7030__S (.I(_3457_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7028__S (.I(_3457_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7141__I0 (.I(_3460_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7122__I0 (.I(_3460_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7054__I0 (.I(_3460_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7033__I0 (.I(_3460_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7143__I0 (.I(_3462_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7124__I0 (.I(_3462_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7056__I0 (.I(_3462_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7036__I0 (.I(_3462_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7246__A2 (.I(_3464_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7227__A2 (.I(_3464_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7187__A2 (.I(_3464_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7039__A1 (.I(_3464_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7056__S (.I(_3465_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7045__I (.I(_3465_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7040__I (.I(_3465_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7053__A2 (.I(_3466_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7052__A2 (.I(_3466_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7043__S (.I(_3466_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7041__S (.I(_3466_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7054__S (.I(_3469_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7050__S (.I(_3469_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7048__S (.I(_3469_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7046__S (.I(_3469_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7116__I (.I(_3500_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7107__I (.I(_3500_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7114__S (.I(_3501_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7112__S (.I(_3501_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7110__S (.I(_3501_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7108__S (.I(_3501_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7124__S (.I(_3506_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7122__S (.I(_3506_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7120__S (.I(_3506_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7117__S (.I(_3506_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7201__I0 (.I(_3508_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7163__I0 (.I(_3508_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7139__I0 (.I(_3508_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7120__I0 (.I(_3508_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7136__I (.I(_3512_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7127__I (.I(_3512_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7134__S (.I(_3513_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7132__S (.I(_3513_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7130__S (.I(_3513_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7128__S (.I(_3513_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7229__I0 (.I(_3523_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7209__I0 (.I(_3523_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7189__I0 (.I(_3523_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7148__I0 (.I(_3523_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7157__S (.I(_3525_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7154__S (.I(_3525_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7151__S (.I(_3525_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7148__S (.I(_3525_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7231__I0 (.I(_3527_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7211__I0 (.I(_3527_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7191__I0 (.I(_3527_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7151__I0 (.I(_3527_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7233__I0 (.I(_3529_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7213__I0 (.I(_3529_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7194__I0 (.I(_3529_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7154__I0 (.I(_3529_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7339__I0 (.I(_3531_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7235__I0 (.I(_3531_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7215__I0 (.I(_3531_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7157__I0 (.I(_3531_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7238__I0 (.I(_3533_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7218__I0 (.I(_3533_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7199__I0 (.I(_3533_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7161__I0 (.I(_3533_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7169__S (.I(_3534_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7166__S (.I(_3534_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7163__S (.I(_3534_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7161__S (.I(_3534_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7242__I0 (.I(_3537_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7223__I0 (.I(_3537_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7203__I0 (.I(_3537_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7166__I0 (.I(_3537_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7244__I0 (.I(_3539_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7225__I0 (.I(_3539_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7205__I0 (.I(_3539_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7169__I0 (.I(_3539_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7198__A2 (.I(_3550_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7197__A2 (.I(_3550_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7191__S (.I(_3550_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7189__S (.I(_3550_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7203__S (.I(_3553_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7201__S (.I(_3553_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7199__S (.I(_3553_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7194__S (.I(_3553_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7318__A1 (.I(_3555_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7295__A1 (.I(_3555_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7254__I1 (.I(_3555_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7197__A1 (.I(_3555_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7217__I (.I(_3561_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7208__I (.I(_3561_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7215__S (.I(_3562_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7213__S (.I(_3562_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7211__S (.I(_3562_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7209__S (.I(_3562_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7225__S (.I(_3567_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7223__S (.I(_3567_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7221__S (.I(_3567_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7218__S (.I(_3567_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7322__I0 (.I(_3569_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7300__I0 (.I(_3569_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7240__I0 (.I(_3569_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7221__I0 (.I(_3569_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7235__S (.I(_3574_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7233__S (.I(_3574_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7231__S (.I(_3574_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7229__S (.I(_3574_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7244__S (.I(_3579_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7242__S (.I(_3579_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7240__S (.I(_3579_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7238__S (.I(_3579_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7256__I (.I(_3584_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7247__I (.I(_3584_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7254__S (.I(_3585_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7252__S (.I(_3585_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7250__S (.I(_3585_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7248__S (.I(_3585_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7263__S (.I(_3590_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7261__S (.I(_3590_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7259__S (.I(_3590_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7257__S (.I(_3590_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7466__I0 (.I(_3603_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7331__I0 (.I(_3603_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7310__I0 (.I(_3603_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7285__I0 (.I(_3603_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7287__I (.I(_3605_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7284__I (.I(_3605_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7298__S (.I(_3606_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7295__A2 (.I(_3606_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7293__A2 (.I(_3606_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7285__S (.I(_3606_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7306__S (.I(_3608_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7303__S (.I(_3608_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7300__S (.I(_3608_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7288__I (.I(_3608_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7597__A1 (.I(_3610_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7554__A1 (.I(_3610_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7314__A1 (.I(_3610_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7290__A1 (.I(_3610_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7599__A1 (.I(_3612_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7556__A1 (.I(_3612_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7316__A1 (.I(_3612_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7293__A1 (.I(_3612_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7476__I0 (.I(_3615_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7342__I0 (.I(_3615_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7320__I0 (.I(_3615_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7298__I0 (.I(_3615_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7480__I0 (.I(_3618_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7347__I0 (.I(_3618_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7324__I0 (.I(_3618_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7303__I0 (.I(_3618_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7482__I0 (.I(_3620_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7349__I0 (.I(_3620_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7326__I0 (.I(_3620_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7306__I0 (.I(_3620_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7312__I (.I(_3622_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7309__I (.I(_3622_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7320__S (.I(_3623_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7318__A2 (.I(_3623_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7316__A2 (.I(_3623_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7310__S (.I(_3623_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7326__S (.I(_3625_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7324__S (.I(_3625_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7322__S (.I(_3625_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7313__I (.I(_3625_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7319__A2 (.I(_3626_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7317__A2 (.I(_3626_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7315__A2 (.I(_3626_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7314__A2 (.I(_3626_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7744__A3 (.I(_3634_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7507__A1 (.I(_3634_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7485__A1 (.I(_3634_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7329__A3 (.I(_3634_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7341__I (.I(_3635_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7330__I (.I(_3635_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7339__S (.I(_3636_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7337__S (.I(_3636_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7334__S (.I(_3636_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7331__S (.I(_3636_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7511__I0 (.I(_3638_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7489__I0 (.I(_3638_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7468__I0 (.I(_3638_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7334__I0 (.I(_3638_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7513__I0 (.I(_3640_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7491__I0 (.I(_3640_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7470__I0 (.I(_3640_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7337__I0 (.I(_3640_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7349__S (.I(_3643_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7347__S (.I(_3643_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7345__S (.I(_3643_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7342__S (.I(_3643_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7520__I0 (.I(_3645_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7499__I0 (.I(_3645_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7478__I0 (.I(_3645_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7345__I0 (.I(_3645_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7763__A2 (.I(_3705_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7570__A1 (.I(_3705_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7526__A2 (.I(_3705_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7464__A2 (.I(_3705_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7473__S (.I(_3707_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7470__S (.I(_3707_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7468__S (.I(_3707_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7466__S (.I(_3707_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7536__I0 (.I(_3711_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7515__I0 (.I(_3711_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7493__I0 (.I(_3711_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7473__I0 (.I(_3711_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7483__I (.I(_3717_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7551__I0 (.I(_3718_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7528__I0 (.I(_3718_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7509__I0 (.I(_3718_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7487__I0 (.I(_3718_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7493__S (.I(_3720_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7491__S (.I(_3720_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7489__S (.I(_3720_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7487__S (.I(_3720_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7561__I0 (.I(_3725_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7539__I0 (.I(_3725_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7518__I0 (.I(_3725_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7497__I0 (.I(_3725_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7505__S (.I(_3726_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7502__S (.I(_3726_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7499__S (.I(_3726_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7497__S (.I(_3726_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7565__I0 (.I(_3729_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7544__I0 (.I(_3729_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7522__I0 (.I(_3729_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7502__I0 (.I(_3729_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7567__I0 (.I(_3731_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7546__I0 (.I(_3731_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7524__I0 (.I(_3731_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7505__I0 (.I(_3731_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7515__S (.I(_3734_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7513__S (.I(_3734_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7511__S (.I(_3734_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7509__S (.I(_3734_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7524__S (.I(_3739_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7522__S (.I(_3739_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7520__S (.I(_3739_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7518__S (.I(_3739_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7536__S (.I(_3745_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7534__S (.I(_3745_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7531__S (.I(_3745_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7528__S (.I(_3745_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7748__I0 (.I(_3747_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7615__I0 (.I(_3747_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7574__I0 (.I(_3747_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7531__I0 (.I(_3747_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7750__I0 (.I(_3749_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7618__I0 (.I(_3749_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7576__I0 (.I(_3749_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7534__I0 (.I(_3749_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7546__S (.I(_3752_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7544__S (.I(_3752_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7542__S (.I(_3752_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7539__S (.I(_3752_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7605__I0 (.I(_3754_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7584__I0 (.I(_3754_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7563__I0 (.I(_3754_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7542__I0 (.I(_3754_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7567__S (.I(_3759_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7565__S (.I(_3759_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7553__I (.I(_3759_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7550__I (.I(_3759_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7563__S (.I(_3760_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7561__S (.I(_3760_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7559__S (.I(_3760_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7551__S (.I(_3760_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7557__A2 (.I(_3762_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7556__A2 (.I(_3762_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7555__A2 (.I(_3762_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7554__A2 (.I(_3762_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7746__I0 (.I(_3771_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7613__I0 (.I(_3771_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7594__I0 (.I(_3771_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7572__I0 (.I(_3771_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7581__I (.I(_3772_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7571__I (.I(_3772_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7578__S (.I(_3773_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7576__S (.I(_3773_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7574__S (.I(_3773_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7572__S (.I(_3773_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7774__I0 (.I(_3778_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7755__I0 (.I(_3778_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7603__I0 (.I(_3778_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7582__I0 (.I(_3778_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7590__S (.I(_3779_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7587__S (.I(_3779_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7584__S (.I(_3779_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7582__S (.I(_3779_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7778__I0 (.I(_3782_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7759__I0 (.I(_3782_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7607__I0 (.I(_3782_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7587__I0 (.I(_3782_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7780__I0 (.I(_3784_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7761__I0 (.I(_3784_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7609__I0 (.I(_3784_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7590__I0 (.I(_3784_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7609__S (.I(_3786_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7607__S (.I(_3786_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7596__I (.I(_3786_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7593__I (.I(_3786_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7605__S (.I(_3787_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7603__S (.I(_3787_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7601__S (.I(_3787_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7594__S (.I(_3787_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7617__I (.I(_3797_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7612__I (.I(_3797_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7630__A2 (.I(_3798_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7628__A2 (.I(_3798_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7615__S (.I(_3798_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7613__S (.I(_3798_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7626__S (.I(_3801_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7622__I (.I(_3801_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7620__S (.I(_3801_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7618__S (.I(_3801_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7795__I0 (.I(_3806_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7776__I0 (.I(_3806_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7757__I0 (.I(_3806_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7626__I0 (.I(_3806_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7754__I (.I(_3866_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7745__I (.I(_3866_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7752__S (.I(_3867_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7750__S (.I(_3867_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7748__S (.I(_3867_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7746__S (.I(_3867_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7771__S (.I(_3878_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7769__S (.I(_3878_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7767__S (.I(_3878_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7765__S (.I(_3878_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7780__S (.I(_3883_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7778__S (.I(_3883_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7776__S (.I(_3883_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7774__S (.I(_3883_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7790__S (.I(_3889_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7788__S (.I(_3889_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7786__S (.I(_3889_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7784__S (.I(_3889_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7829__B (.I(_3908_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7827__A1 (.I(_3908_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7823__A2 (.I(_3908_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7820__A2 (.I(_3908_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7821__I (.I(_3910_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7826__A2 (.I(_3911_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7824__A2 (.I(_3911_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7859__A1 (.I(_3913_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7837__A1 (.I(_3913_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7827__A2 (.I(_3913_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7840__C (.I(_3916_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7835__B (.I(_3916_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7832__I (.I(_3916_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7831__B (.I(_3916_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7861__A1 (.I(_3917_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7860__I (.I(_3917_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7859__A2 (.I(_3917_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7833__A2 (.I(_3917_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1_I (.I(io_in[8]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input2_I (.I(io_in[9]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3987__A2 (.I(\mod.Arithmetic.ACTI.x[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3984__I (.I(\mod.Arithmetic.ACTI.x[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4335__B (.I(\mod.Arithmetic.ACTI.x[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4241__A2 (.I(\mod.Arithmetic.ACTI.x[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4169__A2 (.I(\mod.Arithmetic.ACTI.x[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4071__I (.I(\mod.Arithmetic.ACTI.x[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4453__C (.I(\mod.Arithmetic.ACTI.x[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4336__A2 (.I(\mod.Arithmetic.ACTI.x[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4242__A2 (.I(\mod.Arithmetic.ACTI.x[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4091__I (.I(\mod.Arithmetic.ACTI.x[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4703__C (.I(\mod.Arithmetic.ACTI.x[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4455__A2 (.I(\mod.Arithmetic.ACTI.x[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4104__I (.I(\mod.Arithmetic.ACTI.x[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4767__C (.I(\mod.Arithmetic.ACTI.x[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4704__A2 (.I(\mod.Arithmetic.ACTI.x[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4572__A2 (.I(\mod.Arithmetic.ACTI.x[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4109__I (.I(\mod.Arithmetic.ACTI.x[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4705__A2 (.I(\mod.Arithmetic.ACTI.x[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4597__A1 (.I(\mod.Arithmetic.ACTI.x[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4115__B2 (.I(\mod.Arithmetic.ACTI.x[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4113__B2 (.I(\mod.Arithmetic.ACTI.x[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4768__I0 (.I(\mod.Arithmetic.ACTI.x[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4766__A2 (.I(\mod.Arithmetic.ACTI.x[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4115__A1 (.I(\mod.Arithmetic.ACTI.x[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3996__I (.I(\mod.Arithmetic.ACTI.x[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4038__I (.I(\mod.Arithmetic.CN.I_in[10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4030__I (.I(\mod.Arithmetic.CN.I_in[10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4520__A1 (.I(\mod.Arithmetic.CN.I_in[11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4297__A2 (.I(\mod.Arithmetic.CN.I_in[11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4097__I0 (.I(\mod.Arithmetic.CN.I_in[11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4045__I (.I(\mod.Arithmetic.CN.I_in[11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4517__I (.I(\mod.Arithmetic.CN.I_in[12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4047__I (.I(\mod.Arithmetic.CN.I_in[12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4623__A1 (.I(\mod.Arithmetic.CN.I_in[13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4619__A2 (.I(\mod.Arithmetic.CN.I_in[13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4616__I (.I(\mod.Arithmetic.CN.I_in[13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4054__I (.I(\mod.Arithmetic.CN.I_in[13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4617__I (.I(\mod.Arithmetic.CN.I_in[14] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4060__I (.I(\mod.Arithmetic.CN.I_in[14] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4786__A1 (.I(\mod.Arithmetic.CN.I_in[15] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4067__A1 (.I(\mod.Arithmetic.CN.I_in[15] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3998__I (.I(\mod.Arithmetic.CN.I_in[15] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3967__A2 (.I(\mod.Arithmetic.CN.I_in[16] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3961__I (.I(\mod.Arithmetic.CN.I_in[16] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4127__A2 (.I(\mod.Arithmetic.CN.I_in[17] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4074__I0 (.I(\mod.Arithmetic.CN.I_in[17] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4007__I (.I(\mod.Arithmetic.CN.I_in[17] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4200__A2 (.I(\mod.Arithmetic.CN.I_in[18] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4005__I (.I(\mod.Arithmetic.CN.I_in[18] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4385__A3 (.I(\mod.Arithmetic.CN.I_in[19] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4282__A2 (.I(\mod.Arithmetic.CN.I_in[19] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4003__I (.I(\mod.Arithmetic.CN.I_in[19] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4502__A3 (.I(\mod.Arithmetic.CN.I_in[20] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4501__A2 (.I(\mod.Arithmetic.CN.I_in[20] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4386__A2 (.I(\mod.Arithmetic.CN.I_in[20] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4014__I (.I(\mod.Arithmetic.CN.I_in[20] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4639__A2 (.I(\mod.Arithmetic.CN.I_in[22] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4063__B2 (.I(\mod.Arithmetic.CN.I_in[22] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4018__I (.I(\mod.Arithmetic.CN.I_in[22] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4791__A1 (.I(\mod.Arithmetic.CN.I_in[23] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4025__A1 (.I(\mod.Arithmetic.CN.I_in[23] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4020__A1 (.I(\mod.Arithmetic.CN.I_in[23] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3997__I (.I(\mod.Arithmetic.CN.I_in[23] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4199__A1 (.I(\mod.Arithmetic.CN.I_in[24] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4197__A1 (.I(\mod.Arithmetic.CN.I_in[24] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3969__A2 (.I(\mod.Arithmetic.CN.I_in[24] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3962__A2 (.I(\mod.Arithmetic.CN.I_in[24] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4397__A2 (.I(\mod.Arithmetic.CN.I_in[28] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4389__I (.I(\mod.Arithmetic.CN.I_in[28] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4643__I (.I(\mod.Arithmetic.CN.I_in[30] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4642__A3 (.I(\mod.Arithmetic.CN.I_in[30] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4144__I (.I(\mod.Arithmetic.CN.I_in[32] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3975__A2 (.I(\mod.Arithmetic.CN.I_in[32] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4307__B2 (.I(\mod.Arithmetic.CN.I_in[33] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4153__A3 (.I(\mod.Arithmetic.CN.I_in[33] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4150__A2 (.I(\mod.Arithmetic.CN.I_in[33] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4218__I (.I(\mod.Arithmetic.CN.I_in[34] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4217__A2 (.I(\mod.Arithmetic.CN.I_in[34] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4660__A2 (.I(\mod.Arithmetic.CN.I_in[35] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4543__A1 (.I(\mod.Arithmetic.CN.I_in[35] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4420__A2 (.I(\mod.Arithmetic.CN.I_in[35] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4306__A2 (.I(\mod.Arithmetic.CN.I_in[35] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4542__A2 (.I(\mod.Arithmetic.CN.I_in[36] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4417__I (.I(\mod.Arithmetic.CN.I_in[36] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4755__A1 (.I(\mod.Arithmetic.CN.I_in[37] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4659__I (.I(\mod.Arithmetic.CN.I_in[37] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4632__A1 (.I(\mod.Arithmetic.CN.I_in[37] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4541__A2 (.I(\mod.Arithmetic.CN.I_in[37] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4753__I (.I(\mod.Arithmetic.CN.I_in[38] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4663__A1 (.I(\mod.Arithmetic.CN.I_in[38] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4662__A1 (.I(\mod.Arithmetic.CN.I_in[38] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4756__A1 (.I(\mod.Arithmetic.CN.I_in[39] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4157__A2 (.I(\mod.Arithmetic.CN.I_in[40] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3979__I (.I(\mod.Arithmetic.CN.I_in[40] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4425__A2 (.I(\mod.Arithmetic.CN.I_in[41] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4311__B2 (.I(\mod.Arithmetic.CN.I_in[41] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4157__A3 (.I(\mod.Arithmetic.CN.I_in[41] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4155__A2 (.I(\mod.Arithmetic.CN.I_in[41] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4222__I (.I(\mod.Arithmetic.CN.I_in[42] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4221__A2 (.I(\mod.Arithmetic.CN.I_in[42] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4538__A1 (.I(\mod.Arithmetic.CN.I_in[43] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4309__A2 (.I(\mod.Arithmetic.CN.I_in[43] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4537__A2 (.I(\mod.Arithmetic.CN.I_in[44] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4530__I (.I(\mod.Arithmetic.CN.I_in[44] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4423__A2 (.I(\mod.Arithmetic.CN.I_in[44] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4667__I (.I(\mod.Arithmetic.CN.I_in[45] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4664__A2 (.I(\mod.Arithmetic.CN.I_in[45] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4536__A2 (.I(\mod.Arithmetic.CN.I_in[45] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4751__A2 (.I(\mod.Arithmetic.CN.I_in[46] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4742__A2 (.I(\mod.Arithmetic.CN.I_in[46] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4669__A1 (.I(\mod.Arithmetic.CN.I_in[46] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4665__A1 (.I(\mod.Arithmetic.CN.I_in[46] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4743__A1 (.I(\mod.Arithmetic.CN.I_in[47] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4149__A2 (.I(\mod.Arithmetic.CN.I_in[48] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3981__A2 (.I(\mod.Arithmetic.CN.I_in[48] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4255__I (.I(\mod.Arithmetic.CN.I_in[49] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4162__A2 (.I(\mod.Arithmetic.CN.I_in[49] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4442__A1 (.I(\mod.Arithmetic.CN.I_in[50] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4322__A2 (.I(\mod.Arithmetic.CN.I_in[50] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4253__I (.I(\mod.Arithmetic.CN.I_in[50] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4441__A2 (.I(\mod.Arithmetic.CN.I_in[51] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4323__A2 (.I(\mod.Arithmetic.CN.I_in[51] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4321__A3 (.I(\mod.Arithmetic.CN.I_in[51] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4684__A1 (.I(\mod.Arithmetic.CN.I_in[52] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4553__I (.I(\mod.Arithmetic.CN.I_in[52] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4443__A2 (.I(\mod.Arithmetic.CN.I_in[52] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4440__A1 (.I(\mod.Arithmetic.CN.I_in[52] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4683__I (.I(\mod.Arithmetic.CN.I_in[53] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4557__A1 (.I(\mod.Arithmetic.CN.I_in[53] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4556__A2 (.I(\mod.Arithmetic.CN.I_in[53] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3982__A2 (.I(\mod.Arithmetic.CN.I_in[56] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4439__A2 (.I(\mod.Arithmetic.CN.I_in[57] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4249__A2 (.I(\mod.Arithmetic.CN.I_in[57] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4164__A2 (.I(\mod.Arithmetic.CN.I_in[57] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4555__A2 (.I(\mod.Arithmetic.CN.I_in[58] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4247__I (.I(\mod.Arithmetic.CN.I_in[58] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4555__A3 (.I(\mod.Arithmetic.CN.I_in[59] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4343__I (.I(\mod.Arithmetic.CN.I_in[59] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4769__A3 (.I(\mod.Arithmetic.CN.I_in[61] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4733__A1 (.I(\mod.Arithmetic.CN.I_in[61] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4682__A1 (.I(\mod.Arithmetic.CN.I_in[61] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4578__I (.I(\mod.Arithmetic.CN.I_in[61] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4335__A1 (.I(\mod.Arithmetic.CN.I_in[64] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4234__A3 (.I(\mod.Arithmetic.CN.I_in[64] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3986__A2 (.I(\mod.Arithmetic.CN.I_in[64] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3985__A3 (.I(\mod.Arithmetic.CN.I_in[64] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4703__A1 (.I(\mod.Arithmetic.CN.I_in[67] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4571__A1 (.I(\mod.Arithmetic.CN.I_in[67] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4334__A2 (.I(\mod.Arithmetic.CN.I_in[67] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4767__A1 (.I(\mod.Arithmetic.CN.I_in[68] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4566__A2 (.I(\mod.Arithmetic.CN.I_in[68] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4452__A2 (.I(\mod.Arithmetic.CN.I_in[68] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4746__A1 (.I(\mod.Arithmetic.CN.I_in[69] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4699__A2 (.I(\mod.Arithmetic.CN.I_in[69] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4569__A2 (.I(\mod.Arithmetic.CN.I_in[69] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4749__A2 (.I(\mod.Arithmetic.CN.I_in[70] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4747__I1 (.I(\mod.Arithmetic.CN.I_in[70] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4702__A2 (.I(\mod.Arithmetic.CN.I_in[70] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4745__A2 (.I(\mod.Arithmetic.CN.I_in[71] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4209__A1 (.I(\mod.Arithmetic.CN.I_in[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4208__A1 (.I(\mod.Arithmetic.CN.I_in[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4140__A2 (.I(\mod.Arithmetic.CN.I_in[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3953__I (.I(\mod.Arithmetic.CN.I_in[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4406__A4 (.I(\mod.Arithmetic.CN.I_in[9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4032__I (.I(\mod.Arithmetic.CN.I_in[9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4041__I (.I(\mod.Arithmetic.I_out[72] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4027__I1 (.I(\mod.Arithmetic.I_out[72] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4009__B (.I(\mod.Arithmetic.I_out[72] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4074__I1 (.I(\mod.Arithmetic.I_out[73] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4034__I (.I(\mod.Arithmetic.I_out[73] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4011__B2 (.I(\mod.Arithmetic.I_out[73] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4009__A2 (.I(\mod.Arithmetic.I_out[73] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4031__I1 (.I(\mod.Arithmetic.I_out[74] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4011__A2 (.I(\mod.Arithmetic.I_out[74] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4006__I (.I(\mod.Arithmetic.I_out[74] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6737__I1 (.I(\mod.Data_Mem.F_M.MRAM[0][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6413__I0 (.I(\mod.Data_Mem.F_M.MRAM[0][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6114__B2 (.I(\mod.Data_Mem.F_M.MRAM[0][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6741__I1 (.I(\mod.Data_Mem.F_M.MRAM[0][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6459__A2 (.I(\mod.Data_Mem.F_M.MRAM[0][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5068__I1 (.I(\mod.Data_Mem.F_M.MRAM[0][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6743__I1 (.I(\mod.Data_Mem.F_M.MRAM[0][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6467__A2 (.I(\mod.Data_Mem.F_M.MRAM[0][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5149__I2 (.I(\mod.Data_Mem.F_M.MRAM[0][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6746__I1 (.I(\mod.Data_Mem.F_M.MRAM[0][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6492__A2 (.I(\mod.Data_Mem.F_M.MRAM[0][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5213__I1 (.I(\mod.Data_Mem.F_M.MRAM[0][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6748__I1 (.I(\mod.Data_Mem.F_M.MRAM[0][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6513__A2 (.I(\mod.Data_Mem.F_M.MRAM[0][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5308__A2 (.I(\mod.Data_Mem.F_M.MRAM[0][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6750__I1 (.I(\mod.Data_Mem.F_M.MRAM[0][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6533__A2 (.I(\mod.Data_Mem.F_M.MRAM[0][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5326__I1 (.I(\mod.Data_Mem.F_M.MRAM[0][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6752__I1 (.I(\mod.Data_Mem.F_M.MRAM[0][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6551__A2 (.I(\mod.Data_Mem.F_M.MRAM[0][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5362__I1 (.I(\mod.Data_Mem.F_M.MRAM[0][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7148__I1 (.I(\mod.Data_Mem.F_M.MRAM[12][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6409__A2 (.I(\mod.Data_Mem.F_M.MRAM[12][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6082__B2 (.I(\mod.Data_Mem.F_M.MRAM[12][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7151__I1 (.I(\mod.Data_Mem.F_M.MRAM[12][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6434__A2 (.I(\mod.Data_Mem.F_M.MRAM[12][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6139__B2 (.I(\mod.Data_Mem.F_M.MRAM[12][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7161__I1 (.I(\mod.Data_Mem.F_M.MRAM[12][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6490__I0 (.I(\mod.Data_Mem.F_M.MRAM[12][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6295__B2 (.I(\mod.Data_Mem.F_M.MRAM[12][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7163__I1 (.I(\mod.Data_Mem.F_M.MRAM[12][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6512__A2 (.I(\mod.Data_Mem.F_M.MRAM[12][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6326__B2 (.I(\mod.Data_Mem.F_M.MRAM[12][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7166__I1 (.I(\mod.Data_Mem.F_M.MRAM[12][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6530__A2 (.I(\mod.Data_Mem.F_M.MRAM[12][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6356__B2 (.I(\mod.Data_Mem.F_M.MRAM[12][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7169__I1 (.I(\mod.Data_Mem.F_M.MRAM[12][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6552__A2 (.I(\mod.Data_Mem.F_M.MRAM[12][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6386__B2 (.I(\mod.Data_Mem.F_M.MRAM[12][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6903__I1 (.I(\mod.Data_Mem.F_M.MRAM[13][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6410__A2 (.I(\mod.Data_Mem.F_M.MRAM[13][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6082__A1 (.I(\mod.Data_Mem.F_M.MRAM[13][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6905__I1 (.I(\mod.Data_Mem.F_M.MRAM[13][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6435__A2 (.I(\mod.Data_Mem.F_M.MRAM[13][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6139__A1 (.I(\mod.Data_Mem.F_M.MRAM[13][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6907__I1 (.I(\mod.Data_Mem.F_M.MRAM[13][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6457__A1 (.I(\mod.Data_Mem.F_M.MRAM[13][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6186__A1 (.I(\mod.Data_Mem.F_M.MRAM[13][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6909__I1 (.I(\mod.Data_Mem.F_M.MRAM[13][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6469__A2 (.I(\mod.Data_Mem.F_M.MRAM[13][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6228__A1 (.I(\mod.Data_Mem.F_M.MRAM[13][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6912__I1 (.I(\mod.Data_Mem.F_M.MRAM[13][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6490__I2 (.I(\mod.Data_Mem.F_M.MRAM[13][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6295__A1 (.I(\mod.Data_Mem.F_M.MRAM[13][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6914__I1 (.I(\mod.Data_Mem.F_M.MRAM[13][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6511__A2 (.I(\mod.Data_Mem.F_M.MRAM[13][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6326__A1 (.I(\mod.Data_Mem.F_M.MRAM[13][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6916__I1 (.I(\mod.Data_Mem.F_M.MRAM[13][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6531__A2 (.I(\mod.Data_Mem.F_M.MRAM[13][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6356__A1 (.I(\mod.Data_Mem.F_M.MRAM[13][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6918__I1 (.I(\mod.Data_Mem.F_M.MRAM[13][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6553__A2 (.I(\mod.Data_Mem.F_M.MRAM[13][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6386__A1 (.I(\mod.Data_Mem.F_M.MRAM[13][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6926__I1 (.I(\mod.Data_Mem.F_M.MRAM[14][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6080__A2 (.I(\mod.Data_Mem.F_M.MRAM[14][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5734__I0 (.I(\mod.Data_Mem.F_M.MRAM[14][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6929__I1 (.I(\mod.Data_Mem.F_M.MRAM[14][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6137__A2 (.I(\mod.Data_Mem.F_M.MRAM[14][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5835__I0 (.I(\mod.Data_Mem.F_M.MRAM[14][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6932__I1 (.I(\mod.Data_Mem.F_M.MRAM[14][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6184__A2 (.I(\mod.Data_Mem.F_M.MRAM[14][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5867__I0 (.I(\mod.Data_Mem.F_M.MRAM[14][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6935__I1 (.I(\mod.Data_Mem.F_M.MRAM[14][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6225__A2 (.I(\mod.Data_Mem.F_M.MRAM[14][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5905__I0 (.I(\mod.Data_Mem.F_M.MRAM[14][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6939__I1 (.I(\mod.Data_Mem.F_M.MRAM[14][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6490__I1 (.I(\mod.Data_Mem.F_M.MRAM[14][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6293__B1 (.I(\mod.Data_Mem.F_M.MRAM[14][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5953__A2 (.I(\mod.Data_Mem.F_M.MRAM[14][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6941__I1 (.I(\mod.Data_Mem.F_M.MRAM[14][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6324__B1 (.I(\mod.Data_Mem.F_M.MRAM[14][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5972__I0 (.I(\mod.Data_Mem.F_M.MRAM[14][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6944__I1 (.I(\mod.Data_Mem.F_M.MRAM[14][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6354__B1 (.I(\mod.Data_Mem.F_M.MRAM[14][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6025__I0 (.I(\mod.Data_Mem.F_M.MRAM[14][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6947__I1 (.I(\mod.Data_Mem.F_M.MRAM[14][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6384__B1 (.I(\mod.Data_Mem.F_M.MRAM[14][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6059__I0 (.I(\mod.Data_Mem.F_M.MRAM[14][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6952__I1 (.I(\mod.Data_Mem.F_M.MRAM[15][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6080__B1 (.I(\mod.Data_Mem.F_M.MRAM[15][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5734__I1 (.I(\mod.Data_Mem.F_M.MRAM[15][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4890__A1 (.I(\mod.Data_Mem.F_M.MRAM[15][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6954__I1 (.I(\mod.Data_Mem.F_M.MRAM[15][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6137__B1 (.I(\mod.Data_Mem.F_M.MRAM[15][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5835__I1 (.I(\mod.Data_Mem.F_M.MRAM[15][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4966__B2 (.I(\mod.Data_Mem.F_M.MRAM[15][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6956__I1 (.I(\mod.Data_Mem.F_M.MRAM[15][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6184__B1 (.I(\mod.Data_Mem.F_M.MRAM[15][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5867__I1 (.I(\mod.Data_Mem.F_M.MRAM[15][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5091__B2 (.I(\mod.Data_Mem.F_M.MRAM[15][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6958__I1 (.I(\mod.Data_Mem.F_M.MRAM[15][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6225__B1 (.I(\mod.Data_Mem.F_M.MRAM[15][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5905__I1 (.I(\mod.Data_Mem.F_M.MRAM[15][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5201__A2 (.I(\mod.Data_Mem.F_M.MRAM[15][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6964__I1 (.I(\mod.Data_Mem.F_M.MRAM[15][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6324__A2 (.I(\mod.Data_Mem.F_M.MRAM[15][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5972__I1 (.I(\mod.Data_Mem.F_M.MRAM[15][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5303__A1 (.I(\mod.Data_Mem.F_M.MRAM[15][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6966__I1 (.I(\mod.Data_Mem.F_M.MRAM[15][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6354__A2 (.I(\mod.Data_Mem.F_M.MRAM[15][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6025__I1 (.I(\mod.Data_Mem.F_M.MRAM[15][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5323__A1 (.I(\mod.Data_Mem.F_M.MRAM[15][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6968__I1 (.I(\mod.Data_Mem.F_M.MRAM[15][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6384__A2 (.I(\mod.Data_Mem.F_M.MRAM[15][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6059__I1 (.I(\mod.Data_Mem.F_M.MRAM[15][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5361__A1 (.I(\mod.Data_Mem.F_M.MRAM[15][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6974__I1 (.I(\mod.Data_Mem.F_M.MRAM[16][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5736__I0 (.I(\mod.Data_Mem.F_M.MRAM[16][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4851__I1 (.I(\mod.Data_Mem.F_M.MRAM[16][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6980__I1 (.I(\mod.Data_Mem.F_M.MRAM[16][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5907__I0 (.I(\mod.Data_Mem.F_M.MRAM[16][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5153__I1 (.I(\mod.Data_Mem.F_M.MRAM[16][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6983__I1 (.I(\mod.Data_Mem.F_M.MRAM[16][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5938__I0 (.I(\mod.Data_Mem.F_M.MRAM[16][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5230__I1 (.I(\mod.Data_Mem.F_M.MRAM[16][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6985__I1 (.I(\mod.Data_Mem.F_M.MRAM[16][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5960__I0 (.I(\mod.Data_Mem.F_M.MRAM[16][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5317__I1 (.I(\mod.Data_Mem.F_M.MRAM[16][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6987__I1 (.I(\mod.Data_Mem.F_M.MRAM[16][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6012__I0 (.I(\mod.Data_Mem.F_M.MRAM[16][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5334__I1 (.I(\mod.Data_Mem.F_M.MRAM[16][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6989__I1 (.I(\mod.Data_Mem.F_M.MRAM[16][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6045__I0 (.I(\mod.Data_Mem.F_M.MRAM[16][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5373__I1 (.I(\mod.Data_Mem.F_M.MRAM[16][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6994__I1 (.I(\mod.Data_Mem.F_M.MRAM[17][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5736__I1 (.I(\mod.Data_Mem.F_M.MRAM[17][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4851__I0 (.I(\mod.Data_Mem.F_M.MRAM[17][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6998__I1 (.I(\mod.Data_Mem.F_M.MRAM[17][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5868__I1 (.I(\mod.Data_Mem.F_M.MRAM[17][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5076__I0 (.I(\mod.Data_Mem.F_M.MRAM[17][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7000__I1 (.I(\mod.Data_Mem.F_M.MRAM[17][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5907__I1 (.I(\mod.Data_Mem.F_M.MRAM[17][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5153__I0 (.I(\mod.Data_Mem.F_M.MRAM[17][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7003__I1 (.I(\mod.Data_Mem.F_M.MRAM[17][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5938__I1 (.I(\mod.Data_Mem.F_M.MRAM[17][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5230__I0 (.I(\mod.Data_Mem.F_M.MRAM[17][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7005__I1 (.I(\mod.Data_Mem.F_M.MRAM[17][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5960__I1 (.I(\mod.Data_Mem.F_M.MRAM[17][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5317__I0 (.I(\mod.Data_Mem.F_M.MRAM[17][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7007__I1 (.I(\mod.Data_Mem.F_M.MRAM[17][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6012__I1 (.I(\mod.Data_Mem.F_M.MRAM[17][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5334__I0 (.I(\mod.Data_Mem.F_M.MRAM[17][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7009__I1 (.I(\mod.Data_Mem.F_M.MRAM[17][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6045__I1 (.I(\mod.Data_Mem.F_M.MRAM[17][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5373__I0 (.I(\mod.Data_Mem.F_M.MRAM[17][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7015__I1 (.I(\mod.Data_Mem.F_M.MRAM[18][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5740__I0 (.I(\mod.Data_Mem.F_M.MRAM[18][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4847__I1 (.I(\mod.Data_Mem.F_M.MRAM[18][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7021__I1 (.I(\mod.Data_Mem.F_M.MRAM[18][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5864__I0 (.I(\mod.Data_Mem.F_M.MRAM[18][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5080__I1 (.I(\mod.Data_Mem.F_M.MRAM[18][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7024__I1 (.I(\mod.Data_Mem.F_M.MRAM[18][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5901__I0 (.I(\mod.Data_Mem.F_M.MRAM[18][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5151__I1 (.I(\mod.Data_Mem.F_M.MRAM[18][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7028__I1 (.I(\mod.Data_Mem.F_M.MRAM[18][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5935__I0 (.I(\mod.Data_Mem.F_M.MRAM[18][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5228__I1 (.I(\mod.Data_Mem.F_M.MRAM[18][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7030__I1 (.I(\mod.Data_Mem.F_M.MRAM[18][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5958__I0 (.I(\mod.Data_Mem.F_M.MRAM[18][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5316__I1 (.I(\mod.Data_Mem.F_M.MRAM[18][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7033__I1 (.I(\mod.Data_Mem.F_M.MRAM[18][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6017__A2 (.I(\mod.Data_Mem.F_M.MRAM[18][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5333__I1 (.I(\mod.Data_Mem.F_M.MRAM[18][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7036__I1 (.I(\mod.Data_Mem.F_M.MRAM[18][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6050__A2 (.I(\mod.Data_Mem.F_M.MRAM[18][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5372__I1 (.I(\mod.Data_Mem.F_M.MRAM[18][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7128__I1 (.I(\mod.Data_Mem.F_M.MRAM[19][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5740__I1 (.I(\mod.Data_Mem.F_M.MRAM[19][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4847__I0 (.I(\mod.Data_Mem.F_M.MRAM[19][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7132__I1 (.I(\mod.Data_Mem.F_M.MRAM[19][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5864__I1 (.I(\mod.Data_Mem.F_M.MRAM[19][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5080__I0 (.I(\mod.Data_Mem.F_M.MRAM[19][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7134__I1 (.I(\mod.Data_Mem.F_M.MRAM[19][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5901__I1 (.I(\mod.Data_Mem.F_M.MRAM[19][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5151__I0 (.I(\mod.Data_Mem.F_M.MRAM[19][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7137__I1 (.I(\mod.Data_Mem.F_M.MRAM[19][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5935__I1 (.I(\mod.Data_Mem.F_M.MRAM[19][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5228__I0 (.I(\mod.Data_Mem.F_M.MRAM[19][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7139__I1 (.I(\mod.Data_Mem.F_M.MRAM[19][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5958__I1 (.I(\mod.Data_Mem.F_M.MRAM[19][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5316__I0 (.I(\mod.Data_Mem.F_M.MRAM[19][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7141__I1 (.I(\mod.Data_Mem.F_M.MRAM[19][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6016__A2 (.I(\mod.Data_Mem.F_M.MRAM[19][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5333__I0 (.I(\mod.Data_Mem.F_M.MRAM[19][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7143__I1 (.I(\mod.Data_Mem.F_M.MRAM[19][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6049__A2 (.I(\mod.Data_Mem.F_M.MRAM[19][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5372__I0 (.I(\mod.Data_Mem.F_M.MRAM[19][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7041__I1 (.I(\mod.Data_Mem.F_M.MRAM[1][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6413__I1 (.I(\mod.Data_Mem.F_M.MRAM[1][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6114__A1 (.I(\mod.Data_Mem.F_M.MRAM[1][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7043__I1 (.I(\mod.Data_Mem.F_M.MRAM[1][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6438__I1 (.I(\mod.Data_Mem.F_M.MRAM[1][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4981__I0 (.I(\mod.Data_Mem.F_M.MRAM[1][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7046__I1 (.I(\mod.Data_Mem.F_M.MRAM[1][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6457__B2 (.I(\mod.Data_Mem.F_M.MRAM[1][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5068__I0 (.I(\mod.Data_Mem.F_M.MRAM[1][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7048__I1 (.I(\mod.Data_Mem.F_M.MRAM[1][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6468__A2 (.I(\mod.Data_Mem.F_M.MRAM[1][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6221__I0 (.I(\mod.Data_Mem.F_M.MRAM[1][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5149__I1 (.I(\mod.Data_Mem.F_M.MRAM[1][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7050__I1 (.I(\mod.Data_Mem.F_M.MRAM[1][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6491__A2 (.I(\mod.Data_Mem.F_M.MRAM[1][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5213__I0 (.I(\mod.Data_Mem.F_M.MRAM[1][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7054__I1 (.I(\mod.Data_Mem.F_M.MRAM[1][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6532__A2 (.I(\mod.Data_Mem.F_M.MRAM[1][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5326__I0 (.I(\mod.Data_Mem.F_M.MRAM[1][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7056__I1 (.I(\mod.Data_Mem.F_M.MRAM[1][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6550__A2 (.I(\mod.Data_Mem.F_M.MRAM[1][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5362__I0 (.I(\mod.Data_Mem.F_M.MRAM[1][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7064__I (.I(\mod.Data_Mem.F_M.MRAM[20][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6219__A3 (.I(\mod.Data_Mem.F_M.MRAM[20][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5899__I2 (.I(\mod.Data_Mem.F_M.MRAM[20][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5140__I1 (.I(\mod.Data_Mem.F_M.MRAM[20][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7080__I (.I(\mod.Data_Mem.F_M.MRAM[21][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5899__I3 (.I(\mod.Data_Mem.F_M.MRAM[21][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5140__I0 (.I(\mod.Data_Mem.F_M.MRAM[21][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7175__I (.I(\mod.Data_Mem.F_M.MRAM[22][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6199__A2 (.I(\mod.Data_Mem.F_M.MRAM[22][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5083__A1 (.I(\mod.Data_Mem.F_M.MRAM[22][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7177__I (.I(\mod.Data_Mem.F_M.MRAM[22][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5141__A1 (.I(\mod.Data_Mem.F_M.MRAM[22][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7090__I (.I(\mod.Data_Mem.F_M.MRAM[23][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6119__I0 (.I(\mod.Data_Mem.F_M.MRAM[23][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6692__I1 (.I(\mod.Data_Mem.F_M.MRAM[28][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5665__A2 (.I(\mod.Data_Mem.F_M.MRAM[28][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5567__B2 (.I(\mod.Data_Mem.F_M.MRAM[28][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6696__I1 (.I(\mod.Data_Mem.F_M.MRAM[28][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5673__A2 (.I(\mod.Data_Mem.F_M.MRAM[28][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6701__I1 (.I(\mod.Data_Mem.F_M.MRAM[28][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5688__A2 (.I(\mod.Data_Mem.F_M.MRAM[28][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5595__B2 (.I(\mod.Data_Mem.F_M.MRAM[28][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6705__I1 (.I(\mod.Data_Mem.F_M.MRAM[28][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5699__A2 (.I(\mod.Data_Mem.F_M.MRAM[28][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5604__B2 (.I(\mod.Data_Mem.F_M.MRAM[28][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6709__I1 (.I(\mod.Data_Mem.F_M.MRAM[28][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5709__A2 (.I(\mod.Data_Mem.F_M.MRAM[28][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5611__B2 (.I(\mod.Data_Mem.F_M.MRAM[28][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6713__I1 (.I(\mod.Data_Mem.F_M.MRAM[28][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5720__A2 (.I(\mod.Data_Mem.F_M.MRAM[28][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5618__B2 (.I(\mod.Data_Mem.F_M.MRAM[28][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7189__I1 (.I(\mod.Data_Mem.F_M.MRAM[29][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5632__A2 (.I(\mod.Data_Mem.F_M.MRAM[29][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5524__A1 (.I(\mod.Data_Mem.F_M.MRAM[29][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7191__I1 (.I(\mod.Data_Mem.F_M.MRAM[29][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5650__A2 (.I(\mod.Data_Mem.F_M.MRAM[29][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5552__A1 (.I(\mod.Data_Mem.F_M.MRAM[29][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7194__I1 (.I(\mod.Data_Mem.F_M.MRAM[29][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5663__A2 (.I(\mod.Data_Mem.F_M.MRAM[29][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5567__A1 (.I(\mod.Data_Mem.F_M.MRAM[29][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7199__I1 (.I(\mod.Data_Mem.F_M.MRAM[29][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5685__A2 (.I(\mod.Data_Mem.F_M.MRAM[29][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5595__A1 (.I(\mod.Data_Mem.F_M.MRAM[29][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7201__I1 (.I(\mod.Data_Mem.F_M.MRAM[29][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5697__A2 (.I(\mod.Data_Mem.F_M.MRAM[29][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5604__A1 (.I(\mod.Data_Mem.F_M.MRAM[29][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7203__I1 (.I(\mod.Data_Mem.F_M.MRAM[29][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5708__A2 (.I(\mod.Data_Mem.F_M.MRAM[29][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5611__A1 (.I(\mod.Data_Mem.F_M.MRAM[29][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7205__I1 (.I(\mod.Data_Mem.F_M.MRAM[29][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5718__A2 (.I(\mod.Data_Mem.F_M.MRAM[29][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5618__A1 (.I(\mod.Data_Mem.F_M.MRAM[29][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7209__I1 (.I(\mod.Data_Mem.F_M.MRAM[2][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6112__A2 (.I(\mod.Data_Mem.F_M.MRAM[2][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5743__I0 (.I(\mod.Data_Mem.F_M.MRAM[2][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7211__I1 (.I(\mod.Data_Mem.F_M.MRAM[2][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5827__I0 (.I(\mod.Data_Mem.F_M.MRAM[2][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4980__I1 (.I(\mod.Data_Mem.F_M.MRAM[2][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7213__I1 (.I(\mod.Data_Mem.F_M.MRAM[2][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5863__I0 (.I(\mod.Data_Mem.F_M.MRAM[2][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5072__I1 (.I(\mod.Data_Mem.F_M.MRAM[2][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7218__I1 (.I(\mod.Data_Mem.F_M.MRAM[2][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6493__A2 (.I(\mod.Data_Mem.F_M.MRAM[2][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5949__A2 (.I(\mod.Data_Mem.F_M.MRAM[2][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5215__I1 (.I(\mod.Data_Mem.F_M.MRAM[2][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7221__I1 (.I(\mod.Data_Mem.F_M.MRAM[2][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5971__I0 (.I(\mod.Data_Mem.F_M.MRAM[2][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5310__I1 (.I(\mod.Data_Mem.F_M.MRAM[2][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7223__I1 (.I(\mod.Data_Mem.F_M.MRAM[2][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6024__I0 (.I(\mod.Data_Mem.F_M.MRAM[2][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5327__I1 (.I(\mod.Data_Mem.F_M.MRAM[2][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7225__I1 (.I(\mod.Data_Mem.F_M.MRAM[2][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6055__I0 (.I(\mod.Data_Mem.F_M.MRAM[2][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5364__I1 (.I(\mod.Data_Mem.F_M.MRAM[2][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7229__I1 (.I(\mod.Data_Mem.F_M.MRAM[30][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5522__A2 (.I(\mod.Data_Mem.F_M.MRAM[30][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5463__I0 (.I(\mod.Data_Mem.F_M.MRAM[30][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7231__I1 (.I(\mod.Data_Mem.F_M.MRAM[30][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5834__I0 (.I(\mod.Data_Mem.F_M.MRAM[30][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5550__A2 (.I(\mod.Data_Mem.F_M.MRAM[30][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5473__A2 (.I(\mod.Data_Mem.F_M.MRAM[30][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7235__I1 (.I(\mod.Data_Mem.F_M.MRAM[30][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5580__A2 (.I(\mod.Data_Mem.F_M.MRAM[30][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5481__I0 (.I(\mod.Data_Mem.F_M.MRAM[30][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7238__I1 (.I(\mod.Data_Mem.F_M.MRAM[30][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5593__B1 (.I(\mod.Data_Mem.F_M.MRAM[30][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5492__A2 (.I(\mod.Data_Mem.F_M.MRAM[30][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7240__I1 (.I(\mod.Data_Mem.F_M.MRAM[30][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5602__B1 (.I(\mod.Data_Mem.F_M.MRAM[30][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5499__A2 (.I(\mod.Data_Mem.F_M.MRAM[30][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7242__I1 (.I(\mod.Data_Mem.F_M.MRAM[30][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5609__B1 (.I(\mod.Data_Mem.F_M.MRAM[30][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5505__A2 (.I(\mod.Data_Mem.F_M.MRAM[30][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7244__I1 (.I(\mod.Data_Mem.F_M.MRAM[30][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5616__B1 (.I(\mod.Data_Mem.F_M.MRAM[30][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5512__A2 (.I(\mod.Data_Mem.F_M.MRAM[30][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7248__I0 (.I(\mod.Data_Mem.F_M.MRAM[31][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5522__B1 (.I(\mod.Data_Mem.F_M.MRAM[31][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5463__I1 (.I(\mod.Data_Mem.F_M.MRAM[31][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4890__B1 (.I(\mod.Data_Mem.F_M.MRAM[31][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7252__I0 (.I(\mod.Data_Mem.F_M.MRAM[31][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5565__B1 (.I(\mod.Data_Mem.F_M.MRAM[31][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5477__I1 (.I(\mod.Data_Mem.F_M.MRAM[31][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5091__A2 (.I(\mod.Data_Mem.F_M.MRAM[31][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7257__I0 (.I(\mod.Data_Mem.F_M.MRAM[31][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5593__A2 (.I(\mod.Data_Mem.F_M.MRAM[31][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5491__A2 (.I(\mod.Data_Mem.F_M.MRAM[31][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5222__A1 (.I(\mod.Data_Mem.F_M.MRAM[31][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7259__I0 (.I(\mod.Data_Mem.F_M.MRAM[31][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5602__A2 (.I(\mod.Data_Mem.F_M.MRAM[31][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5501__A2 (.I(\mod.Data_Mem.F_M.MRAM[31][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5313__A1 (.I(\mod.Data_Mem.F_M.MRAM[31][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7261__I0 (.I(\mod.Data_Mem.F_M.MRAM[31][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5609__A2 (.I(\mod.Data_Mem.F_M.MRAM[31][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5504__A2 (.I(\mod.Data_Mem.F_M.MRAM[31][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5330__A1 (.I(\mod.Data_Mem.F_M.MRAM[31][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7263__I0 (.I(\mod.Data_Mem.F_M.MRAM[31][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5616__A2 (.I(\mod.Data_Mem.F_M.MRAM[31][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5511__A2 (.I(\mod.Data_Mem.F_M.MRAM[31][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5369__A1 (.I(\mod.Data_Mem.F_M.MRAM[31][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7108__I1 (.I(\mod.Data_Mem.F_M.MRAM[3][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6113__A2 (.I(\mod.Data_Mem.F_M.MRAM[3][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5743__I1 (.I(\mod.Data_Mem.F_M.MRAM[3][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4876__A1 (.I(\mod.Data_Mem.F_M.MRAM[3][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7112__I1 (.I(\mod.Data_Mem.F_M.MRAM[3][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5863__I1 (.I(\mod.Data_Mem.F_M.MRAM[3][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5072__I0 (.I(\mod.Data_Mem.F_M.MRAM[3][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7114__I1 (.I(\mod.Data_Mem.F_M.MRAM[3][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6221__I2 (.I(\mod.Data_Mem.F_M.MRAM[3][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5902__I1 (.I(\mod.Data_Mem.F_M.MRAM[3][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5149__I0 (.I(\mod.Data_Mem.F_M.MRAM[3][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7117__I1 (.I(\mod.Data_Mem.F_M.MRAM[3][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5948__A2 (.I(\mod.Data_Mem.F_M.MRAM[3][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5215__I0 (.I(\mod.Data_Mem.F_M.MRAM[3][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7120__I1 (.I(\mod.Data_Mem.F_M.MRAM[3][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5971__I1 (.I(\mod.Data_Mem.F_M.MRAM[3][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5310__I0 (.I(\mod.Data_Mem.F_M.MRAM[3][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7122__I1 (.I(\mod.Data_Mem.F_M.MRAM[3][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6024__I1 (.I(\mod.Data_Mem.F_M.MRAM[3][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5327__I0 (.I(\mod.Data_Mem.F_M.MRAM[3][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7124__I1 (.I(\mod.Data_Mem.F_M.MRAM[3][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6055__I1 (.I(\mod.Data_Mem.F_M.MRAM[3][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5364__I0 (.I(\mod.Data_Mem.F_M.MRAM[3][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6881__I (.I(\mod.Data_Mem.F_M.MRAM[4][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5739__I0 (.I(\mod.Data_Mem.F_M.MRAM[4][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4871__I1 (.I(\mod.Data_Mem.F_M.MRAM[4][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6887__I (.I(\mod.Data_Mem.F_M.MRAM[4][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6221__I3 (.I(\mod.Data_Mem.F_M.MRAM[4][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5899__I0 (.I(\mod.Data_Mem.F_M.MRAM[4][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5142__I1 (.I(\mod.Data_Mem.F_M.MRAM[4][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6889__I (.I(\mod.Data_Mem.F_M.MRAM[4][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5950__A2 (.I(\mod.Data_Mem.F_M.MRAM[4][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5209__I1 (.I(\mod.Data_Mem.F_M.MRAM[4][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6891__I (.I(\mod.Data_Mem.F_M.MRAM[4][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5969__A2 (.I(\mod.Data_Mem.F_M.MRAM[4][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5305__I1 (.I(\mod.Data_Mem.F_M.MRAM[4][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6893__I (.I(\mod.Data_Mem.F_M.MRAM[4][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6021__A2 (.I(\mod.Data_Mem.F_M.MRAM[4][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5324__I1 (.I(\mod.Data_Mem.F_M.MRAM[4][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6895__I (.I(\mod.Data_Mem.F_M.MRAM[4][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6057__A2 (.I(\mod.Data_Mem.F_M.MRAM[4][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5365__I1 (.I(\mod.Data_Mem.F_M.MRAM[4][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7271__I (.I(\mod.Data_Mem.F_M.MRAM[5][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5899__I1 (.I(\mod.Data_Mem.F_M.MRAM[5][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5142__I0 (.I(\mod.Data_Mem.F_M.MRAM[5][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7275__I (.I(\mod.Data_Mem.F_M.MRAM[5][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5970__A2 (.I(\mod.Data_Mem.F_M.MRAM[5][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5305__I0 (.I(\mod.Data_Mem.F_M.MRAM[5][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7277__I (.I(\mod.Data_Mem.F_M.MRAM[5][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6022__A2 (.I(\mod.Data_Mem.F_M.MRAM[5][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5324__I0 (.I(\mod.Data_Mem.F_M.MRAM[5][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7279__I (.I(\mod.Data_Mem.F_M.MRAM[5][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6058__A2 (.I(\mod.Data_Mem.F_M.MRAM[5][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5365__I0 (.I(\mod.Data_Mem.F_M.MRAM[5][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6865__I (.I(\mod.Data_Mem.F_M.MRAM[6][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6115__I1 (.I(\mod.Data_Mem.F_M.MRAM[6][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4875__I0 (.I(\mod.Data_Mem.F_M.MRAM[6][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6867__I (.I(\mod.Data_Mem.F_M.MRAM[6][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6144__A2 (.I(\mod.Data_Mem.F_M.MRAM[6][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4975__A1 (.I(\mod.Data_Mem.F_M.MRAM[6][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6869__I (.I(\mod.Data_Mem.F_M.MRAM[6][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6189__A2 (.I(\mod.Data_Mem.F_M.MRAM[6][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5066__A1 (.I(\mod.Data_Mem.F_M.MRAM[6][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7285__I1 (.I(\mod.Data_Mem.F_M.MRAM[768][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5762__A2 (.I(\mod.Data_Mem.F_M.MRAM[768][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4920__I1 (.I(\mod.Data_Mem.F_M.MRAM[768][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7298__I1 (.I(\mod.Data_Mem.F_M.MRAM[768][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6500__A2 (.I(\mod.Data_Mem.F_M.MRAM[768][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5242__I1 (.I(\mod.Data_Mem.F_M.MRAM[768][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7300__I1 (.I(\mod.Data_Mem.F_M.MRAM[768][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6522__A2 (.I(\mod.Data_Mem.F_M.MRAM[768][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5292__A2 (.I(\mod.Data_Mem.F_M.MRAM[768][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7303__I1 (.I(\mod.Data_Mem.F_M.MRAM[768][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6542__A2 (.I(\mod.Data_Mem.F_M.MRAM[768][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5339__I1 (.I(\mod.Data_Mem.F_M.MRAM[768][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7306__I1 (.I(\mod.Data_Mem.F_M.MRAM[768][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6562__A2 (.I(\mod.Data_Mem.F_M.MRAM[768][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5378__I1 (.I(\mod.Data_Mem.F_M.MRAM[768][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6837__I1 (.I(\mod.Data_Mem.F_M.MRAM[769][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6451__A2 (.I(\mod.Data_Mem.F_M.MRAM[769][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5105__A2 (.I(\mod.Data_Mem.F_M.MRAM[769][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6839__I1 (.I(\mod.Data_Mem.F_M.MRAM[769][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6478__A2 (.I(\mod.Data_Mem.F_M.MRAM[769][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5191__A2 (.I(\mod.Data_Mem.F_M.MRAM[769][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6841__I1 (.I(\mod.Data_Mem.F_M.MRAM[769][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6503__A2 (.I(\mod.Data_Mem.F_M.MRAM[769][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5242__I0 (.I(\mod.Data_Mem.F_M.MRAM[769][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6845__I1 (.I(\mod.Data_Mem.F_M.MRAM[769][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6543__A2 (.I(\mod.Data_Mem.F_M.MRAM[769][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5339__I0 (.I(\mod.Data_Mem.F_M.MRAM[769][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6847__I1 (.I(\mod.Data_Mem.F_M.MRAM[769][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6561__B2 (.I(\mod.Data_Mem.F_M.MRAM[769][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5378__I0 (.I(\mod.Data_Mem.F_M.MRAM[769][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7322__I1 (.I(\mod.Data_Mem.F_M.MRAM[770][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5982__I0 (.I(\mod.Data_Mem.F_M.MRAM[770][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5294__I1 (.I(\mod.Data_Mem.F_M.MRAM[770][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7324__I1 (.I(\mod.Data_Mem.F_M.MRAM[770][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6008__I0 (.I(\mod.Data_Mem.F_M.MRAM[770][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5340__I1 (.I(\mod.Data_Mem.F_M.MRAM[770][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7326__I1 (.I(\mod.Data_Mem.F_M.MRAM[770][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6038__I0 (.I(\mod.Data_Mem.F_M.MRAM[770][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5379__I1 (.I(\mod.Data_Mem.F_M.MRAM[770][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7339__I1 (.I(\mod.Data_Mem.F_M.MRAM[771][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5891__A2 (.I(\mod.Data_Mem.F_M.MRAM[771][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5187__A2 (.I(\mod.Data_Mem.F_M.MRAM[771][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7342__I1 (.I(\mod.Data_Mem.F_M.MRAM[771][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5926__I1 (.I(\mod.Data_Mem.F_M.MRAM[771][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5244__I0 (.I(\mod.Data_Mem.F_M.MRAM[771][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7345__I1 (.I(\mod.Data_Mem.F_M.MRAM[771][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5982__I1 (.I(\mod.Data_Mem.F_M.MRAM[771][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5294__I0 (.I(\mod.Data_Mem.F_M.MRAM[771][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7347__I1 (.I(\mod.Data_Mem.F_M.MRAM[771][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6008__I1 (.I(\mod.Data_Mem.F_M.MRAM[771][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5340__I0 (.I(\mod.Data_Mem.F_M.MRAM[771][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7349__I1 (.I(\mod.Data_Mem.F_M.MRAM[771][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6038__I1 (.I(\mod.Data_Mem.F_M.MRAM[771][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5379__I0 (.I(\mod.Data_Mem.F_M.MRAM[771][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7353__I (.I(\mod.Data_Mem.F_M.MRAM[772][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5817__A2 (.I(\mod.Data_Mem.F_M.MRAM[772][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5034__I1 (.I(\mod.Data_Mem.F_M.MRAM[772][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7355__I (.I(\mod.Data_Mem.F_M.MRAM[772][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5856__A2 (.I(\mod.Data_Mem.F_M.MRAM[772][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5095__I1 (.I(\mod.Data_Mem.F_M.MRAM[772][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7369__I (.I(\mod.Data_Mem.F_M.MRAM[773][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5818__A2 (.I(\mod.Data_Mem.F_M.MRAM[773][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5034__I0 (.I(\mod.Data_Mem.F_M.MRAM[773][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7371__I (.I(\mod.Data_Mem.F_M.MRAM[773][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5857__A2 (.I(\mod.Data_Mem.F_M.MRAM[773][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5095__I0 (.I(\mod.Data_Mem.F_M.MRAM[773][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7373__I (.I(\mod.Data_Mem.F_M.MRAM[773][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5893__A2 (.I(\mod.Data_Mem.F_M.MRAM[773][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5182__A2 (.I(\mod.Data_Mem.F_M.MRAM[773][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7405__I (.I(\mod.Data_Mem.F_M.MRAM[775][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5176__A2 (.I(\mod.Data_Mem.F_M.MRAM[775][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7478__I1 (.I(\mod.Data_Mem.F_M.MRAM[780][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6521__A2 (.I(\mod.Data_Mem.F_M.MRAM[780][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6329__B2 (.I(\mod.Data_Mem.F_M.MRAM[780][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7480__I1 (.I(\mod.Data_Mem.F_M.MRAM[780][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6540__A2 (.I(\mod.Data_Mem.F_M.MRAM[780][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6359__B2 (.I(\mod.Data_Mem.F_M.MRAM[780][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7482__I1 (.I(\mod.Data_Mem.F_M.MRAM[780][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6563__A1 (.I(\mod.Data_Mem.F_M.MRAM[780][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6389__B2 (.I(\mod.Data_Mem.F_M.MRAM[780][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7487__I1 (.I(\mod.Data_Mem.F_M.MRAM[781][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6402__A2 (.I(\mod.Data_Mem.F_M.MRAM[781][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6076__A1 (.I(\mod.Data_Mem.F_M.MRAM[781][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7497__I1 (.I(\mod.Data_Mem.F_M.MRAM[781][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6499__I2 (.I(\mod.Data_Mem.F_M.MRAM[781][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6298__A1 (.I(\mod.Data_Mem.F_M.MRAM[781][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7499__I1 (.I(\mod.Data_Mem.F_M.MRAM[781][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6520__A2 (.I(\mod.Data_Mem.F_M.MRAM[781][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6329__A1 (.I(\mod.Data_Mem.F_M.MRAM[781][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7502__I1 (.I(\mod.Data_Mem.F_M.MRAM[781][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6539__A2 (.I(\mod.Data_Mem.F_M.MRAM[781][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6359__A1 (.I(\mod.Data_Mem.F_M.MRAM[781][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7505__I1 (.I(\mod.Data_Mem.F_M.MRAM[781][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6561__A1 (.I(\mod.Data_Mem.F_M.MRAM[781][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6389__A1 (.I(\mod.Data_Mem.F_M.MRAM[781][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7518__I1 (.I(\mod.Data_Mem.F_M.MRAM[782][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6499__I1 (.I(\mod.Data_Mem.F_M.MRAM[782][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6296__B1 (.I(\mod.Data_Mem.F_M.MRAM[782][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5925__I0 (.I(\mod.Data_Mem.F_M.MRAM[782][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7520__I1 (.I(\mod.Data_Mem.F_M.MRAM[782][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6327__B1 (.I(\mod.Data_Mem.F_M.MRAM[782][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5978__A2 (.I(\mod.Data_Mem.F_M.MRAM[782][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7522__I1 (.I(\mod.Data_Mem.F_M.MRAM[782][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6357__B1 (.I(\mod.Data_Mem.F_M.MRAM[782][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6003__A2 (.I(\mod.Data_Mem.F_M.MRAM[782][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7528__I1 (.I(\mod.Data_Mem.F_M.MRAM[783][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6066__B1 (.I(\mod.Data_Mem.F_M.MRAM[783][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5759__I1 (.I(\mod.Data_Mem.F_M.MRAM[783][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4954__B2 (.I(\mod.Data_Mem.F_M.MRAM[783][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7531__I1 (.I(\mod.Data_Mem.F_M.MRAM[783][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6129__A2 (.I(\mod.Data_Mem.F_M.MRAM[783][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5814__I1 (.I(\mod.Data_Mem.F_M.MRAM[783][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5055__A1 (.I(\mod.Data_Mem.F_M.MRAM[783][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7534__I1 (.I(\mod.Data_Mem.F_M.MRAM[783][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6178__A2 (.I(\mod.Data_Mem.F_M.MRAM[783][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5855__I1 (.I(\mod.Data_Mem.F_M.MRAM[783][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5109__A1 (.I(\mod.Data_Mem.F_M.MRAM[783][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7536__I1 (.I(\mod.Data_Mem.F_M.MRAM[783][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6245__A2 (.I(\mod.Data_Mem.F_M.MRAM[783][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5887__A2 (.I(\mod.Data_Mem.F_M.MRAM[783][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5198__A1 (.I(\mod.Data_Mem.F_M.MRAM[783][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7542__I1 (.I(\mod.Data_Mem.F_M.MRAM[783][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6327__A2 (.I(\mod.Data_Mem.F_M.MRAM[783][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5977__A2 (.I(\mod.Data_Mem.F_M.MRAM[783][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5297__A1 (.I(\mod.Data_Mem.F_M.MRAM[783][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7544__I1 (.I(\mod.Data_Mem.F_M.MRAM[783][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6357__A2 (.I(\mod.Data_Mem.F_M.MRAM[783][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6002__A2 (.I(\mod.Data_Mem.F_M.MRAM[783][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5338__A1 (.I(\mod.Data_Mem.F_M.MRAM[783][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7546__I1 (.I(\mod.Data_Mem.F_M.MRAM[783][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6387__A2 (.I(\mod.Data_Mem.F_M.MRAM[783][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6037__I1 (.I(\mod.Data_Mem.F_M.MRAM[783][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5377__A1 (.I(\mod.Data_Mem.F_M.MRAM[783][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7561__I1 (.I(\mod.Data_Mem.F_M.MRAM[784][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5920__I0 (.I(\mod.Data_Mem.F_M.MRAM[784][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5257__I1 (.I(\mod.Data_Mem.F_M.MRAM[784][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7565__I1 (.I(\mod.Data_Mem.F_M.MRAM[784][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5997__I0 (.I(\mod.Data_Mem.F_M.MRAM[784][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5353__I1 (.I(\mod.Data_Mem.F_M.MRAM[784][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7567__I1 (.I(\mod.Data_Mem.F_M.MRAM[784][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6032__I0 (.I(\mod.Data_Mem.F_M.MRAM[784][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5390__I1 (.I(\mod.Data_Mem.F_M.MRAM[784][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7601__I1 (.I(\mod.Data_Mem.F_M.MRAM[786][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5875__I0 (.I(\mod.Data_Mem.F_M.MRAM[786][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5164__I1 (.I(\mod.Data_Mem.F_M.MRAM[786][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7603__I1 (.I(\mod.Data_Mem.F_M.MRAM[786][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5921__A2 (.I(\mod.Data_Mem.F_M.MRAM[786][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5255__A2 (.I(\mod.Data_Mem.F_M.MRAM[786][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7607__I1 (.I(\mod.Data_Mem.F_M.MRAM[786][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5995__A2 (.I(\mod.Data_Mem.F_M.MRAM[786][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5351__A2 (.I(\mod.Data_Mem.F_M.MRAM[786][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7609__I1 (.I(\mod.Data_Mem.F_M.MRAM[786][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6033__A2 (.I(\mod.Data_Mem.F_M.MRAM[786][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5388__A2 (.I(\mod.Data_Mem.F_M.MRAM[786][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7618__I1 (.I(\mod.Data_Mem.F_M.MRAM[787][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5842__A2 (.I(\mod.Data_Mem.F_M.MRAM[787][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5122__A2 (.I(\mod.Data_Mem.F_M.MRAM[787][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7620__I1 (.I(\mod.Data_Mem.F_M.MRAM[787][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5875__I1 (.I(\mod.Data_Mem.F_M.MRAM[787][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5164__I0 (.I(\mod.Data_Mem.F_M.MRAM[787][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7632__I (.I(\mod.Data_Mem.F_M.MRAM[788][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5775__A2 (.I(\mod.Data_Mem.F_M.MRAM[788][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4935__I1 (.I(\mod.Data_Mem.F_M.MRAM[788][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7640__I (.I(\mod.Data_Mem.F_M.MRAM[788][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6283__I3 (.I(\mod.Data_Mem.F_M.MRAM[788][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5917__A2 (.I(\mod.Data_Mem.F_M.MRAM[788][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5251__I1 (.I(\mod.Data_Mem.F_M.MRAM[788][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7646__I (.I(\mod.Data_Mem.F_M.MRAM[788][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6380__I3 (.I(\mod.Data_Mem.F_M.MRAM[788][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6031__A2 (.I(\mod.Data_Mem.F_M.MRAM[788][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5385__I1 (.I(\mod.Data_Mem.F_M.MRAM[788][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6810__I (.I(\mod.Data_Mem.F_M.MRAM[789][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5774__A2 (.I(\mod.Data_Mem.F_M.MRAM[789][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4935__I0 (.I(\mod.Data_Mem.F_M.MRAM[789][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6822__I (.I(\mod.Data_Mem.F_M.MRAM[789][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6341__I0 (.I(\mod.Data_Mem.F_M.MRAM[789][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5993__A2 (.I(\mod.Data_Mem.F_M.MRAM[789][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5347__I2 (.I(\mod.Data_Mem.F_M.MRAM[789][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7648__I (.I(\mod.Data_Mem.F_M.MRAM[790][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6094__A2 (.I(\mod.Data_Mem.F_M.MRAM[790][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4936__A1 (.I(\mod.Data_Mem.F_M.MRAM[790][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7664__I (.I(\mod.Data_Mem.F_M.MRAM[791][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6094__B1 (.I(\mod.Data_Mem.F_M.MRAM[791][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7755__I1 (.I(\mod.Data_Mem.F_M.MRAM[796][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5693__A2 (.I(\mod.Data_Mem.F_M.MRAM[796][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5600__B2 (.I(\mod.Data_Mem.F_M.MRAM[796][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7757__I1 (.I(\mod.Data_Mem.F_M.MRAM[796][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5704__A2 (.I(\mod.Data_Mem.F_M.MRAM[796][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5607__B2 (.I(\mod.Data_Mem.F_M.MRAM[796][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7759__I1 (.I(\mod.Data_Mem.F_M.MRAM[796][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5713__A2 (.I(\mod.Data_Mem.F_M.MRAM[796][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5614__B2 (.I(\mod.Data_Mem.F_M.MRAM[796][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7761__I1 (.I(\mod.Data_Mem.F_M.MRAM[796][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5723__A2 (.I(\mod.Data_Mem.F_M.MRAM[796][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5621__B2 (.I(\mod.Data_Mem.F_M.MRAM[796][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7765__I1 (.I(\mod.Data_Mem.F_M.MRAM[797][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6073__A1 (.I(\mod.Data_Mem.F_M.MRAM[797][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5624__A2 (.I(\mod.Data_Mem.F_M.MRAM[797][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5533__A1 (.I(\mod.Data_Mem.F_M.MRAM[797][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7774__I1 (.I(\mod.Data_Mem.F_M.MRAM[797][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5691__A2 (.I(\mod.Data_Mem.F_M.MRAM[797][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5600__A1 (.I(\mod.Data_Mem.F_M.MRAM[797][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7778__I1 (.I(\mod.Data_Mem.F_M.MRAM[797][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5711__A2 (.I(\mod.Data_Mem.F_M.MRAM[797][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5614__A1 (.I(\mod.Data_Mem.F_M.MRAM[797][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7780__I1 (.I(\mod.Data_Mem.F_M.MRAM[797][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5722__A2 (.I(\mod.Data_Mem.F_M.MRAM[797][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5621__A1 (.I(\mod.Data_Mem.F_M.MRAM[797][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7793__I1 (.I(\mod.Data_Mem.F_M.MRAM[798][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5598__B1 (.I(\mod.Data_Mem.F_M.MRAM[798][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5495__A2 (.I(\mod.Data_Mem.F_M.MRAM[798][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7795__I1 (.I(\mod.Data_Mem.F_M.MRAM[798][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5605__B1 (.I(\mod.Data_Mem.F_M.MRAM[798][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5498__A2 (.I(\mod.Data_Mem.F_M.MRAM[798][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7799__I1 (.I(\mod.Data_Mem.F_M.MRAM[798][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5619__B1 (.I(\mod.Data_Mem.F_M.MRAM[798][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5514__A2 (.I(\mod.Data_Mem.F_M.MRAM[798][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6787__I0 (.I(\mod.Data_Mem.F_M.MRAM[799][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5558__A2 (.I(\mod.Data_Mem.F_M.MRAM[799][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5478__I1 (.I(\mod.Data_Mem.F_M.MRAM[799][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5130__A1 (.I(\mod.Data_Mem.F_M.MRAM[799][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6796__I0 (.I(\mod.Data_Mem.F_M.MRAM[799][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5598__A2 (.I(\mod.Data_Mem.F_M.MRAM[799][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5494__A2 (.I(\mod.Data_Mem.F_M.MRAM[799][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5261__A1 (.I(\mod.Data_Mem.F_M.MRAM[799][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6800__I0 (.I(\mod.Data_Mem.F_M.MRAM[799][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5605__A2 (.I(\mod.Data_Mem.F_M.MRAM[799][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5497__A2 (.I(\mod.Data_Mem.F_M.MRAM[799][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5266__A1 (.I(\mod.Data_Mem.F_M.MRAM[799][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6804__I0 (.I(\mod.Data_Mem.F_M.MRAM[799][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5612__A2 (.I(\mod.Data_Mem.F_M.MRAM[799][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5506__A2 (.I(\mod.Data_Mem.F_M.MRAM[799][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5357__A1 (.I(\mod.Data_Mem.F_M.MRAM[799][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6808__I0 (.I(\mod.Data_Mem.F_M.MRAM[799][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5619__A2 (.I(\mod.Data_Mem.F_M.MRAM[799][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5513__A2 (.I(\mod.Data_Mem.F_M.MRAM[799][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5394__A1 (.I(\mod.Data_Mem.F_M.MRAM[799][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7801__I (.I(\mod.Data_Mem.F_M.MRAM[7][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6115__I0 (.I(\mod.Data_Mem.F_M.MRAM[7][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6922__A1 (.I(\mod.Data_Mem.F_M.dest[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6828__A1 (.I(\mod.Data_Mem.F_M.dest[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6773__A1 (.I(\mod.Data_Mem.F_M.dest[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6677__A1 (.I(\mod.Data_Mem.F_M.dest[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6898__I (.I(\mod.Data_Mem.F_M.dest[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6733__A2 (.I(\mod.Data_Mem.F_M.dest[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6675__A2 (.I(\mod.Data_Mem.F_M.dest[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6970__A1 (.I(\mod.Data_Mem.F_M.dest[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6899__A1 (.I(\mod.Data_Mem.F_M.dest[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6733__A1 (.I(\mod.Data_Mem.F_M.dest[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6675__A1 (.I(\mod.Data_Mem.F_M.dest[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8134__D (.I(\mod.Data_Mem.F_M.out_data[44] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8140__D (.I(\mod.Data_Mem.F_M.out_data[50] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8095__D (.I(\mod.Data_Mem.F_M.out_data[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4872__A1 (.I(\mod.Data_Mem.F_M.src[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4852__I (.I(\mod.Data_Mem.F_M.src[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4833__I (.I(\mod.Data_Mem.F_M.src[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4834__I (.I(\mod.Data_Mem.F_M.src[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4823__I (.I(\mod.Data_Mem.F_M.src[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4885__I (.I(\mod.Data_Mem.F_M.src[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4831__I (.I(\mod.Data_Mem.F_M.src[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4825__I (.I(\mod.Data_Mem.F_M.src[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4865__I (.I(\mod.Data_Mem.F_M.src[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4826__I (.I(\mod.Data_Mem.F_M.src[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5056__I (.I(\mod.Data_Mem.F_M.src[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5001__I (.I(\mod.Data_Mem.F_M.src[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4820__I (.I(\mod.Data_Mem.F_M.src[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7836__A2 (.I(\mod.I_addr[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7819__A2 (.I(\mod.I_addr[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6577__A2 (.I(\mod.I_addr[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6571__I (.I(\mod.I_addr[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4180__A2 (.I(\mod.P2.Rout_reg[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3995__I (.I(\mod.P2.Rout_reg[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3950__A2 (.I(\mod.P2.Rout_reg[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8072__D (.I(\mod.P3.Res[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8073__D (.I(\mod.P3.Res[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8075__D (.I(\mod.P3.Res[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8076__D (.I(\mod.P3.Res[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8077__D (.I(\mod.P3.Res[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8078__D (.I(\mod.P3.Res[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8079__D (.I(\mod.P3.Res[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8595__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8594__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8593__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8592__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8591__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8590__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8589__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8588__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8587__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8586__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8585__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8584__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8583__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8582__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8581__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8580__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8579__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8578__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8577__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8576__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8575__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8574__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8573__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8572__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8571__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8570__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8569__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8568__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8567__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8566__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8565__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8564__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8563__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8562__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8561__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8560__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8559__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8558__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8557__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8556__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8555__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8554__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8553__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8552__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8551__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8550__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8549__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8548__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8547__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8546__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8545__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8544__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8543__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8542__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8541__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8540__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8539__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8538__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8537__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8536__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8535__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8534__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8533__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8532__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8531__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8530__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8529__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8528__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8527__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8526__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8525__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8524__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8523__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8522__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8521__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8520__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8519__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8518__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8517__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8516__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8515__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8514__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8513__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8512__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8511__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8510__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8509__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8508__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8507__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8506__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8505__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8504__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8503__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8502__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8501__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8500__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8499__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8498__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8497__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8496__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8495__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8494__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8493__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8492__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8491__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8490__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8489__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8488__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8487__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8486__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8485__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8484__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8483__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8482__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8481__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8480__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8479__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8478__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8477__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8476__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8475__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8474__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8473__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8472__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8471__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8470__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8469__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8468__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8467__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8466__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8465__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8464__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8463__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8462__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8461__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8460__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8459__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8458__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8457__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8456__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8455__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8454__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8453__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8452__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8451__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8450__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8449__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8448__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8447__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8446__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8445__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8444__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8443__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8442__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8441__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8440__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8439__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8438__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8437__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8436__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8435__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8434__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8433__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8432__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8431__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8430__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8429__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8428__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8427__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8426__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8425__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8424__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8423__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8422__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8421__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8420__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8419__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8418__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8417__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8416__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8415__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8414__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8413__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8412__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8411__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8410__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8409__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8408__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8407__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8406__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8405__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8404__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8403__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8402__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8401__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8400__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8399__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8398__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8397__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8396__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8395__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8394__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8393__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8392__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8391__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8390__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8389__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8388__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8387__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8386__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8385__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8384__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8383__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8382__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8381__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8380__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8379__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8378__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8377__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8376__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8375__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8374__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8373__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8372__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8371__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8370__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8369__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8368__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8367__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8366__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8365__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8364__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8363__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8362__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8361__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8360__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8359__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8358__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8357__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8356__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8355__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8354__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8353__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8352__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8351__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8350__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8349__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8348__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8347__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8346__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8345__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8344__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8343__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8342__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8341__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8340__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8339__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8338__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8337__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8336__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8335__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8334__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8333__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8332__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8331__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8330__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8329__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8328__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8327__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8326__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8325__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8324__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8323__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8322__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8321__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8320__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8319__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8318__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8317__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8316__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8315__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8314__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8313__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8312__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8311__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8310__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8309__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8308__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8307__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8306__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8305__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8304__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8303__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8302__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8301__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8300__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8299__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8298__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8297__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8296__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8295__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8294__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8293__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8292__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8291__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8290__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8289__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8288__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8287__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8286__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8285__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8284__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8283__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8282__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8281__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8280__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8279__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8278__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8277__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8276__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8275__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8274__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8273__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8272__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8271__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8270__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8269__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8268__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8267__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8266__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8265__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8264__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8263__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8262__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8261__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8260__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8259__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8258__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8257__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8256__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8255__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8254__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8253__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8252__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8251__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8250__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8249__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8248__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8247__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8246__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8245__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8244__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8243__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8242__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8241__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8240__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8239__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8238__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8237__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8236__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8235__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8234__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8233__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8232__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8231__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8230__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8229__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8228__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8227__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8226__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8225__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8224__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8223__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8222__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8221__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8220__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8219__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8218__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8217__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8216__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8215__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8214__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8213__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8212__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8211__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8210__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8209__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8208__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8207__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8206__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8205__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8204__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8203__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8202__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8201__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8200__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8199__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8198__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8197__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8196__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8195__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8194__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8193__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8192__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8191__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8190__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8189__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8188__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8187__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8186__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8185__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8184__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8183__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8182__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8181__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8180__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8179__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8178__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8177__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8176__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8175__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8174__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8173__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8172__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8171__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8170__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8169__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8168__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8167__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8166__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8165__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8164__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8163__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8162__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8161__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8160__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8159__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8158__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8157__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8156__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8155__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8154__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8153__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8152__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8151__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8150__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8149__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8148__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8147__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8146__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8145__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8144__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8143__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8142__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8141__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8140__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8139__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8138__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8137__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8136__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8135__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8134__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8133__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8132__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8131__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8130__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8129__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8128__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8127__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8126__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8125__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8124__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8123__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8122__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8121__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8120__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8119__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8118__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8117__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8116__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8115__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8114__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8113__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8112__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8111__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8110__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8109__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8108__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8107__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8106__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8105__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8104__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8103__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8102__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8101__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8100__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8099__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8098__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8097__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8096__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8095__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8094__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8093__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8092__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8091__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8090__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8089__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8088__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8087__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8086__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8085__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8084__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8083__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8082__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8081__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8080__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8079__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8078__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8077__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8076__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8075__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8074__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8073__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8072__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8071__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8070__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8069__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8068__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8067__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8066__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8065__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8064__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8063__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8062__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8061__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8060__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8059__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8058__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8057__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8056__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8055__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8054__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8053__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8052__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8051__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8050__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8049__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8048__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8047__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8046__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8045__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8044__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8043__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8042__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8041__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8040__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8039__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8038__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8037__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8036__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8035__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8034__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8033__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8032__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8031__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8030__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8029__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8028__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8027__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8026__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8025__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8024__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8023__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8022__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8021__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8020__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8019__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8018__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8017__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8016__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8015__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8014__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8013__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8012__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8011__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8010__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8009__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8008__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8007__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8006__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8005__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8004__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8003__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8002__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8001__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8000__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7999__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7998__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7997__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7996__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7995__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7994__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7993__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7992__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7991__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7990__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7989__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7988__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7987__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7986__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7985__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7984__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7983__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7982__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7981__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7980__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7979__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7978__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7977__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7976__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7975__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7974__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7973__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7972__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7971__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7970__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7969__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7968__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7967__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7966__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7965__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7964__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7963__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7962__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7961__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7960__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7959__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7958__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7957__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7956__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7955__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7954__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7953__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7952__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7951__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7950__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7949__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7948__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7947__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7946__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7945__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7944__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7943__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7942__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7941__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7940__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7939__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7938__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7937__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7936__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7935__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7934__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7933__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7932__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7931__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7930__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7929__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7928__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7927__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7926__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7925__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7924__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7923__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7922__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7921__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7920__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7919__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7918__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7917__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7916__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7915__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7914__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7913__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7912__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7911__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7910__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7909__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7908__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7907__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7906__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7905__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7904__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7903__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7902__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7901__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7900__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7899__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7898__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7897__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7896__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7895__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7894__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7893__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7892__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7891__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7890__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7889__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7888__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7887__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7886__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7885__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7884__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7883__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7882__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7881__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7880__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7879__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7878__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7877__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7876__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7875__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7874__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7873__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7872__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7871__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7870__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7869__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7868__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7867__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7866__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7865__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7864__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7863__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7862__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8231__RN (.I(net2));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8230__RN (.I(net2));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8229__RN (.I(net2));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8228__RN (.I(net2));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8227__RN (.I(net2));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8202__RN (.I(net2));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8201__RN (.I(net2));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8200__RN (.I(net2));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8199__RN (.I(net2));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8198__RN (.I(net2));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8197__RN (.I(net2));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8196__RN (.I(net2));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8195__RN (.I(net2));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8194__RN (.I(net2));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8177__RN (.I(net2));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8176__RN (.I(net2));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8175__RN (.I(net2));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8174__RN (.I(net2));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8173__RN (.I(net2));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8172__RN (.I(net2));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8171__RN (.I(net2));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8170__RN (.I(net2));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8169__RN (.I(net2));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8168__RN (.I(net2));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8167__RN (.I(net2));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8166__RN (.I(net2));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8165__RN (.I(net2));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8164__RN (.I(net2));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8163__RN (.I(net2));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8162__RN (.I(net2));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8161__RN (.I(net2));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8160__RN (.I(net2));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8159__RN (.I(net2));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8158__RN (.I(net2));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8157__RN (.I(net2));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8156__RN (.I(net2));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8155__RN (.I(net2));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8154__RN (.I(net2));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8153__RN (.I(net2));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8152__RN (.I(net2));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8151__RN (.I(net2));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8150__RN (.I(net2));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8149__RN (.I(net2));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8148__RN (.I(net2));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8147__RN (.I(net2));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8146__RN (.I(net2));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8145__RN (.I(net2));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8144__RN (.I(net2));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8143__RN (.I(net2));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8142__RN (.I(net2));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8141__RN (.I(net2));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8140__RN (.I(net2));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8139__RN (.I(net2));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8138__RN (.I(net2));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8137__RN (.I(net2));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8136__RN (.I(net2));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8135__RN (.I(net2));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8134__RN (.I(net2));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8133__RN (.I(net2));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8132__RN (.I(net2));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8131__RN (.I(net2));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8130__RN (.I(net2));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8129__RN (.I(net2));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8128__RN (.I(net2));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8127__RN (.I(net2));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8126__RN (.I(net2));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8125__RN (.I(net2));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8124__RN (.I(net2));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8123__RN (.I(net2));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8122__RN (.I(net2));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8121__RN (.I(net2));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8120__RN (.I(net2));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8119__RN (.I(net2));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8118__RN (.I(net2));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8117__RN (.I(net2));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8116__RN (.I(net2));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8115__RN (.I(net2));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8114__RN (.I(net2));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8113__RN (.I(net2));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8112__RN (.I(net2));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8111__RN (.I(net2));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8110__RN (.I(net2));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8109__RN (.I(net2));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8108__RN (.I(net2));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8107__RN (.I(net2));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8106__RN (.I(net2));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8105__RN (.I(net2));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8104__RN (.I(net2));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8103__RN (.I(net2));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8102__RN (.I(net2));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8101__RN (.I(net2));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8100__RN (.I(net2));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8099__RN (.I(net2));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8098__RN (.I(net2));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8097__RN (.I(net2));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8096__RN (.I(net2));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8095__RN (.I(net2));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8094__RN (.I(net2));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8093__RN (.I(net2));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8092__RN (.I(net2));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8091__RN (.I(net2));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8090__RN (.I(net2));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8089__RN (.I(net2));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8088__RN (.I(net2));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8079__RN (.I(net2));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8078__RN (.I(net2));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8077__RN (.I(net2));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8076__RN (.I(net2));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8075__RN (.I(net2));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8074__RN (.I(net2));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8073__RN (.I(net2));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8072__RN (.I(net2));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8071__RN (.I(net2));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7998__RN (.I(net2));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7997__RN (.I(net2));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7996__RN (.I(net2));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7995__RN (.I(net2));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7994__RN (.I(net2));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7993__RN (.I(net2));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7992__RN (.I(net2));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7991__RN (.I(net2));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7990__RN (.I(net2));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7989__RN (.I(net2));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7988__RN (.I(net2));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7987__RN (.I(net2));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7986__RN (.I(net2));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7985__RN (.I(net2));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7984__RN (.I(net2));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7983__RN (.I(net2));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7982__RN (.I(net2));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output3_I (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6770__I (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6673__I (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output4_I (.I(net4));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6781__I (.I(net4));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6686__I (.I(net4));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output5_I (.I(net5));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6785__I (.I(net5));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6690__I (.I(net5));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output6_I (.I(net6));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6789__I (.I(net6));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6694__I (.I(net6));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output7_I (.I(net7));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6793__I (.I(net7));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6698__I (.I(net7));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output8_I (.I(net8));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6798__I (.I(net8));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6703__I (.I(net8));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output9_I (.I(net9));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6802__I (.I(net9));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6707__I (.I(net9));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output10_I (.I(net10));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6806__I (.I(net10));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6711__I (.I(net10));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_17 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_77 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_145 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_287 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_462 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_497 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_533 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_569 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_678 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1073 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_1092 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1127 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1172 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1178 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_1_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_462 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_1_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_1_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_1_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_2_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_2_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_2_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_2_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_497 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_2_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_2_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_2_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_2_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_3_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_3_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_3_532 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_3_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_4_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_4_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_4_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_4_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_4_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_4_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_4_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_4_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_4_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_5_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_5_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_5_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_6_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_6_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_6_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_6_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_6_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_6_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_6_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_6_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_7_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_8_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_8_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_8_571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_8_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_8_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_1213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_9_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_9_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_9_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_9_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_10_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_10_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_10_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_568 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_571 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_10_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_10_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_10_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_1213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_11_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_11_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_11_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_11_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_11_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_11_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_12_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_12_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_12_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_12_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_355 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_429 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_12_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_1207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_13_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_13_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_603 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_607 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_610 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_13_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_13_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_14_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_14_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_429 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_14_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_14_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_14_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_14_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_14_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_14_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_14_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_15_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_15_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_572 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_610 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_15_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_15_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_15_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_15_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_15_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_15_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_16_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_429 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_498 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_16_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_16_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_16_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_17_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_17_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_433 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_674 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_17_678 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_17_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_17_751 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_17_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_17_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_18_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_18_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_18_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_18_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_571 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_643 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_18_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_18_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_18_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_19_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_319 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_674 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_678 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_19_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_19_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_19_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_20_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_20_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_20_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_20_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_639 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_643 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_678 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_20_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_20_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_20_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_1213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_319 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_21_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_21_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_21_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_22_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_22_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_22_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_22_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_569 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_607 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_642 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_22_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_22_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_22_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_1213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_23_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_23_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_320 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_464 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_643 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_23_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_23_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_24_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_285 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_571 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_24_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_24_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_24_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_25_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_25_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_461 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_607 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_25_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_25_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_26_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_26_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_26_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_26_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_497 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_568 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_713 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_26_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_26_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_27_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_461 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_606 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_27_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_27_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_28_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_28_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_28_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_28_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_320 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_532 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_29_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_29_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_29_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_30_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_30_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_30_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_285 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_642 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_30_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_822 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_30_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_30_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_30_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_30_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_31_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_31_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_533 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_31_752 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_31_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_31_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_32_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_32_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_32_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_355 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_32_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_32_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_32_878 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_32_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_32_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_33_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_33_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_33_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_390 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_33_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_33_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_33_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_33_913 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_33_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_34_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_34_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_427 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_498 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_571 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_642 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_34_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_34_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_34_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_34_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_34_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_810 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_34_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_1085 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_34_1089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_34_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_34_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_35_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_35_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_249 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_606 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_610 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_35_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_678 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_748 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_35_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_35_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_36_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_36_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_36_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_36_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_36_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_36_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_1035 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_1080 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_36_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_36_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_1207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_532 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_603 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_607 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_37_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_37_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_748 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_37_752 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_37_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_37_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_38_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_38_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_287 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_427 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_569 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_38_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_713 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_38_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_38_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_38_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_852 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_38_855 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_38_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_923 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_38_926 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_38_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_38_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_39_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_39_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_604 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_39_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_39_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_674 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_677 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_39_890 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_39_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_39_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_39_964 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_39_980 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_39_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_40_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_642 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_40_713 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_40_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_40_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_40_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_40_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_878 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_924 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_40_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_40_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_987 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_995 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_40_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_40_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_40_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_40_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_41_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_248 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_390 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_533 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_41_610 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_41_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_678 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_41_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_748 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_752 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_41_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_41_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_806 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_41_810 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_41_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_41_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_41_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_878 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_890 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_964 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_981 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_985 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_41_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_41_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_1059 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_41_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_42_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_42_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_42_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_42_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_42_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_42_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_42_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_569 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_42_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_42_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_42_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_703 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_805 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_42_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_42_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_42_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_875 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_878 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_980 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_984 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_1000 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_1016 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_1020 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_42_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_42_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_1213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_43_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_43_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_43_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_43_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_249 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_319 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_464 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_604 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_674 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_43_678 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_43_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_43_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_806 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_810 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_816 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_43_819 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_43_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_843 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_915 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_981 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_985 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_1035 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_43_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_43_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_43_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_44_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_44_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_44_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_44_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_429 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_568 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_44_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_44_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_44_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_44_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_987 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_995 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_44_1050 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_44_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_44_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_44_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_45_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_45_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_45_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_45_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_462 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_45_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_45_610 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_45_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_45_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_45_806 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_816 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_964 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_972 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_974 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_981 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_985 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1053 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1057 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_45_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_46_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_46_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_46_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_46_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_46_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_46_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_46_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_46_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_46_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_572 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_46_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_678 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_711 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_46_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_46_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_46_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_822 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_845 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_972 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_983 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_987 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1066 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_46_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_46_1090 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_46_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_46_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_46_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_1213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_47_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_390 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_47_394 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_47_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_461 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_47_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_47_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_47_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_47_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_47_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_47_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_47_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_604 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_606 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_47_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_47_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_677 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_47_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_703 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_47_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_47_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_751 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_47_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_817 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_820 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_910 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_962 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1050 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_47_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_47_1110 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_47_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_47_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_48_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_48_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_48_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_48_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_48_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_48_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_213 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_48_285 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_427 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_48_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_48_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_497 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_48_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_48_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_703 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_751 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_48_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_855 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_946 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_950 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_994 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1059 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1075 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_48_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_48_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_48_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_48_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_1213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_49_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_49_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_49_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_49_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_49_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_322 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_49_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_49_464 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_49_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_49_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_49_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_572 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_603 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_49_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_49_738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_746 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_805 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_816 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_910 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_964 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_981 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_985 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1029 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1051 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1090 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_49_1094 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_49_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_49_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_50_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_50_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_50_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_50_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_50_285 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_50_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_50_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_50_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_429 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_50_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_50_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_50_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_50_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_703 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_50_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_50_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_781 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_891 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_894 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_910 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_913 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_981 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_985 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1050 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1068 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1072 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1080 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1088 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1092 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_50_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_50_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_50_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_51_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_51_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_248 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_51_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_51_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_462 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_51_533 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_572 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_603 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_607 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_51_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_51_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_703 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_51_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_51_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_816 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_820 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_864 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_911 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_981 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_985 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_1050 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_1090 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_1094 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_51_1110 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_51_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_51_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_52_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_52_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_52_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_52_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_52_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_285 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_52_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_52_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_52_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_52_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_52_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_569 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_52_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_52_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_52_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_639 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_642 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_52_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_678 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_52_713 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_52_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_52_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_822 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_929 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1050 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_1068 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_1072 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1090 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1094 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_52_1121 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_52_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_52_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_52_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_53_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_53_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_53_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_53_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_249 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_53_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_53_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_53_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_53_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_53_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_53_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_53_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_53_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_53_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_53_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_603 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_53_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_643 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_53_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_53_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_820 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_911 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_915 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_964 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_974 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_1029 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_1053 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_1085 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_1089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_1093 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_1123 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_53_1127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_53_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_53_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_54_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_54_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_54_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_54_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_54_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_54_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_54_571 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_54_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_54_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_54_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_54_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_781 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_54_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_924 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_1107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_54_1140 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_54_1156 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_1164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_54_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_54_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_55_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_55_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_55_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_55_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_462 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_55_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_55_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_55_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_55_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_606 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_55_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_55_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_677 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_55_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_748 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_55_752 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_55_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_55_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_819 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_867 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_959 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_987 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_1020 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_1030 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_1032 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_1058 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_1073 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_1093 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_1104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_1108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_55_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_55_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_55_1193 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_1201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_55_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_56_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_56_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_56_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_56_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_56_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_56_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_429 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_497 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_56_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_568 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_56_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_56_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_56_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_56_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_56_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_56_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_56_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_822 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_878 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_985 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_1000 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_1053 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_1055 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_1094 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_1137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_56_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_56_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_56_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_57_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_57_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_248 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_57_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_57_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_57_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_57_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_461 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_532 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_604 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_57_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_57_677 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_746 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_810 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_984 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_1018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_1051 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_1058 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_1108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_1123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_1127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_57_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_57_1197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_57_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_58_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_58_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_58_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_217 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_287 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_58_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_569 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_820 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_924 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_945 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_981 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_985 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1000 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1020 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1055 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1066 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_1080 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_58_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_58_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_1213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_59_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_59_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_83 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_59_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_59_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_533 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_607 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_59_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_59_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_59_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_703 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_59_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_59_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_817 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_891 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_945 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_962 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_974 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_984 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1030 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1057 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_1101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_1110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_1114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_59_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_59_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_60_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_60_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_60_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_60_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_60_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_60_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_60_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_60_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_60_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_60_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_60_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_60_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_643 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_678 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_60_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_60_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_840 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_962 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_995 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1020 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_60_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_60_1208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_61_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_61_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_61_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_319 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_61_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_61_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_464 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_61_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_61_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_61_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_61_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_61_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_61_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_61_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_61_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_61_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_745 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_819 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1016 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1080 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1090 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_1104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_1125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1195 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_61_1199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_61_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_62_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_62_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_62_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_62_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_62_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_62_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_607 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_610 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_62_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_62_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_713 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_62_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_62_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_781 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_806 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_820 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_891 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_910 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_927 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_948 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1016 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1050 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1069 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_1073 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_1085 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_62_1208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_17 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_63_21 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_63_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_63_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_249 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_63_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_63_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_461 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_464 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_63_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_533 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_63_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_674 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_677 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_703 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_63_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_745 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_748 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_816 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_820 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_891 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_930 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_985 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1080 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_1094 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_63_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_64_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_64_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_64_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_77 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_64_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_64_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_429 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_64_433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_64_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_64_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_568 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_571 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_64_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_64_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_806 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_820 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_913 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_929 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_945 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_965 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1020 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1050 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1069 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_1104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_1167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_65_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_65_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_319 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_65_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_65_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_65_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_65_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_532 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_65_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_65_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_65_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_65_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_65_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_65_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_751 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_816 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_822 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_830 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_891 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_894 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_910 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_931 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_950 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_964 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1030 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1058 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1080 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1094 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_1104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1128 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_66_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_66_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_66_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_285 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_355 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_359 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_66_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_66_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_427 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_66_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_66_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_497 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_66_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_66_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_568 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_66_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_639 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_711 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_66_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_66_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_782 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_820 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_878 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_891 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_910 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_974 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_987 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_995 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1057 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1072 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_67_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_67_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_87 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_178 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_248 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_67_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_67_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_67_461 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_67_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_67_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_703 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_67_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_748 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_67_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_819 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_959 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_965 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_1016 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1032 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1085 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_68_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_68_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_71 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_74 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_217 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_68_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_427 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_68_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_68_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_68_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_568 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_678 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_68_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_68_713 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_68_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_751 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_68_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_782 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_840 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_894 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_911 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_924 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_1018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1085 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_69_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_69_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_69_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_462 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_69_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_532 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_603 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_607 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_69_677 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_69_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_806 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_810 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_820 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_894 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_911 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_930 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_961 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1090 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_1092 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_1203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_70_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_70_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_70_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_70_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_70_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_70_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_70_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_70_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_70_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_70_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_642 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_70_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_703 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_70_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_70_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_70_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_878 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_910 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_931 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_997 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1072 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1092 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_71_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_71_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_71_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_71_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_71_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_572 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_71_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_71_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_819 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_911 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_985 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1030 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_1032 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1053 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1094 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_1110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_1203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_72_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_72_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_72_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_72_429 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_72_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_569 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_642 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_72_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_782 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_810 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_891 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_945 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_962 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_974 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_984 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_1000 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1050 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1075 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1090 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_73_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_73_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_73_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_73_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_533 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_603 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_607 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_610 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_73_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_73_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_73_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_73_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_843 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_946 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_972 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_1020 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_1050 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1094 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1178 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_74_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_74_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_74_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_74_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_429 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_497 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_607 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_610 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_74_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_74_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_751 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_805 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_822 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_830 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_878 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_880 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_894 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_910 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_926 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_945 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_994 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1093 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1160 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_1167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_75_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_75_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_75_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_75_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_178 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_75_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_319 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_75_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_75_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_532 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_674 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_678 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_75_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_75_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_746 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_817 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_891 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_980 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1059 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_76_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_76_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_76_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_76_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_76_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_76_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_76_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_497 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_607 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_639 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_76_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_678 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_751 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_945 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_983 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1016 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1058 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1075 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_77_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_77_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_77_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_77_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_77_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_77_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_77_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_77_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_77_462 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_77_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_77_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_748 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_817 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_946 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_965 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_981 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_985 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1032 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1055 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1178 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_78_5 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_78_21 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_29 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_78_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_214 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_78_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_78_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_78_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_497 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_639 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_643 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_78_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_78_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_782 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_878 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_880 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_924 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_985 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_997 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_1057 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1068 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1080 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1094 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_1123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1210 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_1214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_79_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_79_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_79_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_79_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_532 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_603 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_606 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_610 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_79_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_79_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_806 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_810 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_864 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_911 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_945 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_984 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1020 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1032 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_1051 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_1055 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_80_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_80_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_80_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_80_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_80_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_80_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_80_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_948 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_998 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1059 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_1127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1211 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_1215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_81_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_81_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_81_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_81_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_81_462 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_81_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_572 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_604 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_745 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_751 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_845 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_915 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_984 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1050 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_82_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_82_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_82_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_82_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_82_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_82_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_711 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_820 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_891 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_894 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_930 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_945 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_985 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1050 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_1085 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_1167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_83_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_83_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_83_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_83_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_572 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_703 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_746 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_819 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_915 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1020 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1059 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_1093 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_1203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_84_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_84_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_84_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_427 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_429 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_639 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_713 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_84_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_810 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_830 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_867 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_878 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_894 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_985 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_995 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_997 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1069 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1094 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_1167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_85_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_85_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_85_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_85_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_85_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_320 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_604 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_607 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_85_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_677 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_85_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_745 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_85_748 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_806 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_819 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_843 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_915 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1058 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1090 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_1123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1178 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_86_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_86_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_86_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_86_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_86_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_284 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_427 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_497 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_86_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_643 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_711 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_713 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_852 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_855 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_903 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_995 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1055 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1072 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_87_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_87_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_87_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_87_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_87_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_87_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_87_322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_603 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_643 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_87_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_87_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_87_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_87_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_87_748 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_806 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_819 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_915 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1016 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1029 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1178 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_88_5 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_88_21 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_29 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_88_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_88_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_88_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_88_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_88_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_287 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_88_291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_88_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_355 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_88_568 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_88_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_88_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_88_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_88_713 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_88_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_88_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_782 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_843 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1050 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1066 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_1075 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_88_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_89_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_89_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_89_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_89_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_89_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_462 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_464 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_89_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_89_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_89_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_746 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_820 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_1029 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1055 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1080 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_1088 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_89_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_90_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_90_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_90_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_90_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_90_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_90_213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_90_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_90_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_90_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_90_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_90_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_355 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_90_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_90_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_643 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_90_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_90_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_90_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_781 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_806 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_867 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_878 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_962 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_981 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_995 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1051 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1071 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_1073 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_1104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1196 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_90_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_90_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_91_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_91_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_91_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_91_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_91_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_249 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_91_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_91_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_320 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_91_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_91_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_91_603 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_91_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_91_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_677 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_91_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_745 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_91_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_816 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_820 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_867 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_913 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_915 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_984 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_1051 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_91_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_91_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_92_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_92_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_92_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_355 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_569 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_643 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_92_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_92_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_711 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_713 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_92_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_92_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_92_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_92_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_830 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_876 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_880 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_1066 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1093 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_92_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_92_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_93_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_93_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_93_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_93_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_93_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_93_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_249 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_320 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_674 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_93_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_93_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_93_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_751 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_93_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_845 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_930 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1029 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1058 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1075 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1090 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_1100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_93_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_1201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_93_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_94_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_94_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_94_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_94_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_285 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_94_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_568 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_572 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_639 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_643 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_806 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_852 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_856 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1057 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1066 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_94_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_94_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_94_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_95_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_95_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_95_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_95_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_95_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_95_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_95_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_461 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_572 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_678 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_745 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_820 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_984 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1030 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_1090 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_95_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_95_1181 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_95_1197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_95_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_96_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_96_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_96_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_96_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_96_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_96_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_355 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_96_359 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_96_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_96_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_96_433 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_569 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_96_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_782 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_931 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_1020 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1085 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_96_1139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_96_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_96_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_1213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_97_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_97_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_97_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_97_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_97_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_249 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_97_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_97_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_319 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_97_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_390 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_97_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_462 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_97_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_677 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_97_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_97_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_746 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_806 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_810 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_817 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_819 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_987 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1093 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_97_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_97_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_98_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_98_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_98_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_217 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_98_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_284 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_98_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_98_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_711 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_782 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_98_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_810 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_845 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_945 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_995 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_997 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1020 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1093 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1121 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_98_1125 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_98_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_98_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_98_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_99_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_99_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_99_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_99_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_99_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_248 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_359 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_533 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_607 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_99_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_674 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_748 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_99_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_99_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_99_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_810 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_819 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_948 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1059 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1114 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_99_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_99_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_99_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_100_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_100_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_100_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_100_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_100_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_284 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_100_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_100_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_100_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_355 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_569 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_100_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_100_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_100_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_100_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_100_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_782 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_100_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_806 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_875 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_878 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_924 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_962 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1077 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1088 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1092 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_100_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_100_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_100_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_100_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_100_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_101_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_101_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_101_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_101_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_101_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_101_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_101_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_101_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_101_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_101_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_532 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_610 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_674 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_101_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_101_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_101_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_101_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_101_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_101_819 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_101_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_913 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_915 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_981 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1055 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1080 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1094 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_101_1110 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_101_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_101_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_101_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_102_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_102_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_102_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_214 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_102_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_102_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_102_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_102_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_571 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_102_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_102_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_102_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_102_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_102_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_751 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_781 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_102_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_830 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_102_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_995 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1090 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1094 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_102_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_102_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_102_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_1213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_103_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_103_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_103_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_103_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_103_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_103_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_464 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_674 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_678 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_703 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_103_746 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_822 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_103_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_103_888 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_910 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_930 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_987 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1088 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1092 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_103_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_103_1128 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_103_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_103_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_104_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_104_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_104_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_104_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_104_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_285 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_427 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_610 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_104_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_855 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_104_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_867 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_104_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_104_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_104_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_913 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_915 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_964 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1000 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1051 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1055 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_104_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_104_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_104_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_105_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_105_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_105_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_105_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_105_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_319 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_390 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_533 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_105_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_105_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_105_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_105_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_105_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_105_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_105_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_105_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_915 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1055 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1059 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_105_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_1129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_105_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_105_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_106_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_106_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_106_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_106_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_284 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_106_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_427 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_498 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_569 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_639 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_642 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_678 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_106_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_106_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_106_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_106_805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_106_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_106_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_106_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_913 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_948 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_965 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_972 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_1051 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_106_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_1094 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_106_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_106_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_106_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_107_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_107_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_107_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_107_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_107_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_107_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_107_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_107_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_107_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_107_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_107_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_959 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_981 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_985 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1050 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1058 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_107_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_107_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_107_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_107_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_107_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_108_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_108_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_108_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_108_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_285 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_429 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_713 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_108_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_108_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_108_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_806 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_108_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_108_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_867 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_108_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_913 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_948 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_108_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_987 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_994 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_998 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_108_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1020 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_108_1065 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_108_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_108_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_108_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_1213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_109_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_109_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_109_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_109_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_109_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_249 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_572 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_606 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_746 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_109_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_109_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_843 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_109_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_109_974 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_109_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1032 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_109_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_109_1050 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_1058 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_109_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_109_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_109_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_110_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_110_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_110_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_110_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_355 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_497 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_782 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_110_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_110_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_110_931 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_110_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_110_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_110_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_110_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_110_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_110_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_111_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_111_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_111_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_111_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_532 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_604 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_607 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_111_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_748 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_111_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_111_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_111_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_810 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_816 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_111_819 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_843 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_111_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_111_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_111_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_927 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_111_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_111_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_111_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_111_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_111_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_111_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_112_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_112_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_112_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_568 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_643 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_112_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_112_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_112_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_112_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_880 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_112_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_112_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_964 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_995 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_112_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_112_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_112_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_112_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_112_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_112_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_113_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_113_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_113_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_113_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_113_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_533 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_677 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_113_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_113_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_113_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_113_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_113_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_113_984 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_998 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_113_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_113_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_113_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_113_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_113_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_17 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_114_21 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_29 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_114_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_114_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_114_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_114_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_427 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_711 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_114_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_114_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_114_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_114_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_820 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_114_843 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_114_875 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_114_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_114_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_948 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_950 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_114_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_114_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_114_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_1093 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_114_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_114_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_114_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_115_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_115_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_115_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_610 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_678 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_115_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_115_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_115_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_115_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_115_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_115_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_115_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_115_983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_115_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_115_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_115_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_1058 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_115_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_115_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_115_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_116_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_116_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_116_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_429 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_498 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_568 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_116_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_116_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_116_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_116_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_116_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_931 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_116_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_116_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_116_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_116_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_116_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_116_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_117_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_117_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_117_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_117_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_117_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_117_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_572 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_606 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_117_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_117_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_751 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_117_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_117_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_117_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_816 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_820 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_117_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_117_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_117_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_894 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_117_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_117_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_117_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_117_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_985 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_117_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_117_1035 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_117_1051 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_1059 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_117_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_117_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_117_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_118_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_118_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_118_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_118_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_355 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_118_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_118_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_118_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_118_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_118_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_118_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_118_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_118_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_118_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_911 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_915 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_118_950 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_118_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_974 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_118_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_118_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_118_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_118_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_118_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_118_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_1213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_119_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_119_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_119_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_119_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_119_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_461 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_572 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_119_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_119_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_119_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_119_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_888 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_891 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_119_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_119_945 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_119_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_985 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_119_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_119_1035 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_119_1051 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_1059 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_119_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_119_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_119_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_120_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_120_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_120_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_120_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_120_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_120_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_429 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_498 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_120_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_120_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_751 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_120_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_120_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_120_806 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_120_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_120_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_120_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_120_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_120_948 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_120_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_974 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_120_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_120_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_120_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_120_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_120_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_120_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_1213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_121_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_121_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_121_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_121_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_121_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_121_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_572 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_121_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_121_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_121_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_822 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_121_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_843 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_121_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_864 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_121_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_121_911 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_121_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_121_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_121_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_121_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_121_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_122_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_122_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_122_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_122_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_122_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_122_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_122_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_122_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_569 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_122_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_122_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_122_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_122_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_122_856 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_122_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_880 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_122_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_122_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_122_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_122_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_122_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_122_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_122_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_122_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_123_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_123_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_123_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_123_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_123_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_123_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_123_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_123_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_123_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_123_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_390 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_607 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_123_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_123_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_830 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_123_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_123_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_123_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_123_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_123_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_987 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_123_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_123_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_123_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_123_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_124_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_124_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_124_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_124_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_124_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_124_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_607 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_610 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_124_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_124_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_124_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_124_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_124_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_124_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_124_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_124_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_124_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_124_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_124_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_124_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_124_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_124_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_125_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_125_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_125_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_125_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_125_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_125_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_125_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_125_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_390 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_606 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_610 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_125_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_125_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_125_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_125_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_805 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_125_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_125_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_125_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_125_911 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_125_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_125_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_125_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_125_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_125_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_126_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_126_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_126_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_126_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_126_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_126_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_355 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_126_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_126_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_126_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_751 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_126_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_126_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_126_806 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_126_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_875 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_126_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_126_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_948 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_126_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_126_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_127_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_127_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_127_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_127_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_127_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_461 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_127_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_127_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_127_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_127_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_127_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_127_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_127_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_127_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_127_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_127_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_127_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_127_843 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_127_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_127_915 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_127_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_127_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_127_983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_127_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_128_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_128_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_128_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_128_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_77 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_128_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_128_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_118 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_128_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_128_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_128_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_128_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_128_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_128_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_429 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_569 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_128_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_128_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_128_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_128_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_128_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_128_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_128_864 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_880 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_128_926 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_128_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_128_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_128_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_128_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_128_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_1213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_129_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_129_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_129_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_129_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_129_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_129_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_129_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_129_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_129_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_129_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_129_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_129_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_129_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_129_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_129_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_129_604 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_129_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_129_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_129_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_845 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_129_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_129_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_878 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_129_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_129_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_910 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_129_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_130_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_130_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_130_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_130_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_130_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_130_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_130_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_130_359 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_130_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_130_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_130_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_130_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_130_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_130_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_130_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_130_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_130_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_130_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_130_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_130_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_130_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_810 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_130_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_852 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_855 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_130_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_130_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_130_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_130_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_130_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_130_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_131_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_131_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_249 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_131_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_319 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_131_322 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_131_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_131_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_131_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_131_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_131_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_131_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_131_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_131_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_131_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_131_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_131_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_131_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_131_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_131_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_131_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_131_913 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_929 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_131_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_131_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_987 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_131_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_132_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_132_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_132_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_132_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_132_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_132_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_132_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_132_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_132_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_132_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_132_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_132_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_132_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_132_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_751 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_132_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_132_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_132_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_132_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_132_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_132_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_132_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_974 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_132_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_132_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_132_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_132_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_133_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_133_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_133_55 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_133_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_133_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_133_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_133_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_133_249 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_133_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_133_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_133_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_133_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_133_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_133_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_133_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_133_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_133_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_133_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_133_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_748 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_133_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_133_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_133_830 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_133_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_891 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_133_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_948 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_133_964 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_133_980 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_133_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_133_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_133_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_134_40 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_48 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_52 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_134_83 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_134_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_134_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_134_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_134_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_134_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_134_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_134_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_134_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_134_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_134_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_134_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_134_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_134_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_134_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_134_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_134_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_134_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_134_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_134_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_134_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_134_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_134_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_134_806 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_134_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_134_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_134_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_915 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_134_923 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_134_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_134_1000 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_134_1016 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_134_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_134_1071 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_134_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_134_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_134_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_135_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_135_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_135_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_135_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_135_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_135_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_135_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_135_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_135_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_135_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_135_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_135_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_135_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_135_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_806 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_810 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_817 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_135_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_135_880 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_890 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_135_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_135_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_135_1050 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_1058 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_135_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_136_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_136_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_136_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_77 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_136_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_136_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_136_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_136_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_136_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_136_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_136_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_136_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_136_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_903 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_136_910 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_136_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_136_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_136_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_77 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_79 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_82 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_137_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_137_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_137_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_138_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_138_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_138_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_1213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_139_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_140_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_140_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_140_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_1213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_141_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_142_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_142_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_142_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_142_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_143_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_144_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_144_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_144_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_144_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_144_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_144_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_144_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_144_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_144_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_144_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_144_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_144_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_144_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_144_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_144_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_144_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_144_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_144_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_1207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_145_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_145_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_145_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_145_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_145_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_145_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_145_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_145_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_145_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_145_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_145_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_145_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_145_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_145_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_145_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_145_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_145_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_145_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_145_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_145_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_145_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_145_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_145_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_145_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_145_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_145_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_145_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_145_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_145_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_145_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_145_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_145_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_145_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_145_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_145_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_145_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_146_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_146_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_146_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_146_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_146_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_146_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_146_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_146_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_146_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_146_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_146_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_146_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_146_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_146_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_146_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_146_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_146_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_146_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_146_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_147_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_147_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_147_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_147_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_147_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_147_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_147_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_147_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_147_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_147_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_147_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_147_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_147_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_147_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_147_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_147_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_147_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_147_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_148_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_148_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_148_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_148_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_148_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_148_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_148_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_148_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_148_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_148_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_148_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_148_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_148_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_148_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_148_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_148_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_148_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_148_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_148_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_149_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_149_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_149_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_149_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_149_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_149_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_149_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_149_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_149_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_149_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_149_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_149_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_149_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_149_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_149_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_149_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_149_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_149_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_149_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_149_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_149_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_149_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_149_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_149_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_149_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_149_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_149_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_149_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_149_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_149_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_149_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_149_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_149_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_149_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_149_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_150_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_150_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_150_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_150_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_150_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_150_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_150_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_150_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_150_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_150_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_150_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_150_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_150_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_150_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_150_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_150_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_150_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_150_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_150_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_150_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_151_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_151_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_151_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_151_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_151_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_151_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_151_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_151_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_151_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_151_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_151_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_151_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_151_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_151_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_151_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_151_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_151_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_151_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_151_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_151_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_151_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_151_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_151_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_151_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_151_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_151_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_151_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_151_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_151_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_151_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_151_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_151_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_151_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_151_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_151_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_151_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_152_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_152_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_152_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_152_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_152_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_152_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_152_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_152_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_152_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_152_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_152_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_152_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_152_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_152_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_152_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_152_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_152_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_152_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_152_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_152_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_152_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_152_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_152_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_152_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_152_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_152_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_152_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_152_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_152_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_152_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_152_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_152_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_152_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_152_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_152_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_153_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_153_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_153_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_153_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_153_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_153_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_153_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_153_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_153_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_153_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_153_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_153_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_153_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_153_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_153_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_153_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_153_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_153_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_153_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_153_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_153_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_153_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_153_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_153_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_153_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_153_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_153_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_153_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_153_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_153_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_153_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_153_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_153_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_153_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_153_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_153_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_154_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_154_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_154_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_154_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_154_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_154_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_154_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_154_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_154_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_154_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_154_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_154_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_154_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_154_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_154_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_154_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_154_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_154_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_154_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_154_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_154_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_154_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_154_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_154_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_154_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_154_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_154_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_154_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_154_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_154_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_154_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_154_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_154_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_154_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_154_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_155_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_155_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_155_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_155_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_155_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_155_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_155_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_155_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_155_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_155_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_155_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_155_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_155_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_155_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_155_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_155_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_155_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_155_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_156_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_156_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_156_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_156_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_156_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_156_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_156_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_156_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_156_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_156_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_156_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_156_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_156_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_156_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_156_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_156_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_156_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_156_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_156_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_156_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_156_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_156_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_156_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_156_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_156_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_156_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_156_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_156_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_156_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_156_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_156_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_156_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_156_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_156_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_156_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_157_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_157_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_157_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_157_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_157_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_157_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_157_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_157_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_157_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_157_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_157_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_157_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_157_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_157_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_157_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_157_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_157_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_157_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_158_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_158_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_158_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_158_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_158_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_158_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_158_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_158_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_158_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_158_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_158_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_158_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_158_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_158_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_158_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_158_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_158_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_158_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_158_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_158_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_158_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_158_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_158_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_158_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_158_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_158_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_158_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_158_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_158_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_158_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_158_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_158_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_158_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_158_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_158_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_159_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_159_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_159_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_159_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_159_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_159_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_159_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_159_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_159_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_159_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_159_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_159_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_159_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_159_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_159_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_159_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_159_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_159_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_159_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_159_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_159_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_159_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_159_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_159_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_159_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_159_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_159_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_159_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_159_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_159_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_159_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_159_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_159_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_159_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_159_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_159_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_160_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_160_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_160_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_160_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_160_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_160_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_160_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_160_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_160_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_160_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_160_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_160_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_160_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_160_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_160_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_160_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_160_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_160_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_160_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_160_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_160_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_160_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_160_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_160_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_160_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_160_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_160_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_160_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_160_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_160_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_160_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_160_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_160_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_160_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_160_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_160_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_161_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_161_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_161_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_161_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_161_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_161_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_161_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_161_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_161_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_161_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_161_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_161_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_161_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_161_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_161_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_161_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_161_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_161_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_161_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_161_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_161_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_161_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_161_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_161_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_161_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_161_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_161_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_161_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_161_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_161_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_161_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_161_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_161_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_161_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_161_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_161_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_162_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_162_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_162_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_162_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_162_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_162_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_162_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_162_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_162_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_162_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_162_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_162_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_162_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_162_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_162_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_162_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_162_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_162_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_162_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_162_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_162_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_162_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_162_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_162_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_162_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_162_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_162_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_162_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_162_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_162_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_162_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_162_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_162_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_162_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_162_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_162_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_163_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_163_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_163_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_163_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_163_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_163_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_163_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_163_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_163_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_163_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_163_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_163_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_163_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_163_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_163_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_163_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_163_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_163_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_163_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_163_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_163_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_163_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_163_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_163_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_163_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_163_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_163_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_163_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_163_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_163_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_163_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_163_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_163_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_163_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_163_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_163_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_163_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_164_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_164_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_164_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_164_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_164_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_164_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_164_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_164_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_164_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_164_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_164_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_164_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_164_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_164_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_164_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_164_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_164_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_164_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_164_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_165_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_165_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_165_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_165_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_165_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_165_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_165_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_165_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_165_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_165_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_165_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_165_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_165_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_165_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_165_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_165_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_165_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_165_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_165_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_165_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_165_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_165_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_165_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_165_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_165_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_165_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_165_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_165_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_165_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_165_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_165_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_165_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_165_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_165_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_165_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_165_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_165_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_165_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_165_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_165_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_165_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_165_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_165_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_165_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_165_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_165_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_165_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_165_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_165_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_165_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_165_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_165_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_165_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_165_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_165_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_166_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_166_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_166_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_166_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_166_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_166_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_166_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_166_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_166_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_166_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_166_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_166_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_166_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_166_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_166_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_166_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_166_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_166_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_166_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_166_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_166_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_166_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_166_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_166_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_166_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_166_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_166_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_166_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_166_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_166_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_166_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_166_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_166_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_166_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_166_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_166_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_166_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_166_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_167_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_167_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_167_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_167_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_167_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_167_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_167_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_167_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_167_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_167_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_167_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_167_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_167_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_167_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_167_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_167_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_167_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_167_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_167_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_167_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_167_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_167_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_167_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_167_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_167_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_167_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_167_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_167_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_167_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_167_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_167_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_167_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_167_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_167_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_167_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_167_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_167_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_167_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_167_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_167_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_167_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_167_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_167_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_167_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_167_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_167_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_167_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_167_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_167_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_167_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_167_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_167_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_167_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_167_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_167_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_168_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_168_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_168_13 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_168_29 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_168_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_168_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_168_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_168_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_168_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_168_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_168_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_168_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_168_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_168_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_168_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_168_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_168_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_168_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_168_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_168_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_168_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_168_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_168_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_168_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_168_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_168_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_168_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_168_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_168_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_168_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_168_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_168_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_168_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_168_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_168_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_168_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_168_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_168_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_168_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_168_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_168_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_168_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_168_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_168_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_168_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_168_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_168_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_168_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_168_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_168_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_168_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_168_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_168_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_168_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_168_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_168_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_168_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_169_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_169_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_169_11 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_169_17 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_169_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_169_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_169_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_169_42 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_169_46 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_169_48 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_169_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_169_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_169_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_169_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_169_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_169_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_169_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_169_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_169_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_169_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_169_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_169_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_169_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_169_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_169_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_169_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_169_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_169_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_169_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_169_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_169_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_169_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_169_285 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_169_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_169_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_169_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_169_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_169_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_169_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_169_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_169_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_169_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_169_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_169_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_169_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_169_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_169_427 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_169_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_169_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_169_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_169_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_169_462 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_169_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_169_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_169_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_169_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_169_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_169_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_169_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_169_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_169_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_169_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_169_569 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_169_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_169_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_169_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_169_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_169_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_169_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_169_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_169_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_169_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_169_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_169_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_169_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_169_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_169_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_169_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_169_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_169_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_169_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_169_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_169_713 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_169_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_169_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_169_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_169_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_169_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_169_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_169_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_169_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_169_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_169_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_169_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_169_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_169_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_169_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_169_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_169_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_169_852 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_169_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_169_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_169_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_169_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_169_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_169_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_169_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_169_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_169_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_169_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_169_924 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_169_929 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_169_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_169_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_169_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_169_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_169_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_169_994 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_169_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_169_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_169_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_169_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_169_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_169_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_169_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_169_1068 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_169_1073 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_169_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_169_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_169_1092 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_169_1108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_169_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_169_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_169_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_169_1128 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_169_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_169_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_169_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_169_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_169_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_169_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_169_1197 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_169_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_169_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_169_1223 ();
 assign io_oeb[0] = net11;
 assign io_oeb[10] = net21;
 assign io_oeb[11] = net22;
 assign io_oeb[12] = net23;
 assign io_oeb[13] = net24;
 assign io_oeb[14] = net25;
 assign io_oeb[15] = net26;
 assign io_oeb[16] = net27;
 assign io_oeb[17] = net28;
 assign io_oeb[18] = net29;
 assign io_oeb[19] = net30;
 assign io_oeb[1] = net12;
 assign io_oeb[20] = net31;
 assign io_oeb[21] = net32;
 assign io_oeb[22] = net33;
 assign io_oeb[23] = net34;
 assign io_oeb[24] = net35;
 assign io_oeb[25] = net36;
 assign io_oeb[26] = net37;
 assign io_oeb[27] = net38;
 assign io_oeb[28] = net39;
 assign io_oeb[29] = net40;
 assign io_oeb[2] = net13;
 assign io_oeb[30] = net41;
 assign io_oeb[31] = net42;
 assign io_oeb[32] = net43;
 assign io_oeb[33] = net44;
 assign io_oeb[34] = net45;
 assign io_oeb[35] = net46;
 assign io_oeb[36] = net47;
 assign io_oeb[37] = net48;
 assign io_oeb[3] = net14;
 assign io_oeb[4] = net15;
 assign io_oeb[5] = net16;
 assign io_oeb[6] = net17;
 assign io_oeb[7] = net18;
 assign io_oeb[8] = net19;
 assign io_oeb[9] = net20;
 assign io_out[0] = net49;
 assign io_out[10] = net59;
 assign io_out[11] = net60;
 assign io_out[12] = net61;
 assign io_out[13] = net62;
 assign io_out[14] = net63;
 assign io_out[15] = net64;
 assign io_out[1] = net50;
 assign io_out[24] = net65;
 assign io_out[25] = net66;
 assign io_out[26] = net67;
 assign io_out[27] = net68;
 assign io_out[28] = net69;
 assign io_out[29] = net70;
 assign io_out[2] = net51;
 assign io_out[30] = net71;
 assign io_out[31] = net72;
 assign io_out[32] = net73;
 assign io_out[33] = net74;
 assign io_out[34] = net75;
 assign io_out[35] = net76;
 assign io_out[36] = net77;
 assign io_out[37] = net78;
 assign io_out[3] = net52;
 assign io_out[4] = net53;
 assign io_out[5] = net54;
 assign io_out[6] = net55;
 assign io_out[7] = net56;
 assign io_out[8] = net57;
 assign io_out[9] = net58;
 assign la_data_out[0] = net79;
 assign la_data_out[10] = net89;
 assign la_data_out[11] = net90;
 assign la_data_out[12] = net91;
 assign la_data_out[13] = net92;
 assign la_data_out[14] = net93;
 assign la_data_out[15] = net94;
 assign la_data_out[16] = net95;
 assign la_data_out[17] = net96;
 assign la_data_out[18] = net97;
 assign la_data_out[19] = net98;
 assign la_data_out[1] = net80;
 assign la_data_out[20] = net99;
 assign la_data_out[21] = net100;
 assign la_data_out[22] = net101;
 assign la_data_out[23] = net102;
 assign la_data_out[24] = net103;
 assign la_data_out[25] = net104;
 assign la_data_out[26] = net105;
 assign la_data_out[27] = net106;
 assign la_data_out[28] = net107;
 assign la_data_out[29] = net108;
 assign la_data_out[2] = net81;
 assign la_data_out[30] = net109;
 assign la_data_out[31] = net110;
 assign la_data_out[32] = net111;
 assign la_data_out[33] = net112;
 assign la_data_out[34] = net113;
 assign la_data_out[35] = net114;
 assign la_data_out[36] = net115;
 assign la_data_out[37] = net116;
 assign la_data_out[38] = net117;
 assign la_data_out[39] = net118;
 assign la_data_out[3] = net82;
 assign la_data_out[40] = net119;
 assign la_data_out[41] = net120;
 assign la_data_out[42] = net121;
 assign la_data_out[43] = net122;
 assign la_data_out[44] = net123;
 assign la_data_out[45] = net124;
 assign la_data_out[46] = net125;
 assign la_data_out[47] = net126;
 assign la_data_out[48] = net127;
 assign la_data_out[49] = net128;
 assign la_data_out[4] = net83;
 assign la_data_out[50] = net129;
 assign la_data_out[51] = net130;
 assign la_data_out[52] = net131;
 assign la_data_out[53] = net132;
 assign la_data_out[54] = net133;
 assign la_data_out[55] = net134;
 assign la_data_out[56] = net135;
 assign la_data_out[57] = net136;
 assign la_data_out[58] = net137;
 assign la_data_out[59] = net138;
 assign la_data_out[5] = net84;
 assign la_data_out[60] = net139;
 assign la_data_out[61] = net140;
 assign la_data_out[62] = net141;
 assign la_data_out[63] = net142;
 assign la_data_out[6] = net85;
 assign la_data_out[7] = net86;
 assign la_data_out[8] = net87;
 assign la_data_out[9] = net88;
 assign user_irq[0] = net143;
 assign user_irq[1] = net144;
 assign user_irq[2] = net145;
 assign wbs_ack_o = net146;
 assign wbs_dat_o[0] = net147;
 assign wbs_dat_o[10] = net157;
 assign wbs_dat_o[11] = net158;
 assign wbs_dat_o[12] = net159;
 assign wbs_dat_o[13] = net160;
 assign wbs_dat_o[14] = net161;
 assign wbs_dat_o[15] = net162;
 assign wbs_dat_o[16] = net163;
 assign wbs_dat_o[17] = net164;
 assign wbs_dat_o[18] = net165;
 assign wbs_dat_o[19] = net166;
 assign wbs_dat_o[1] = net148;
 assign wbs_dat_o[20] = net167;
 assign wbs_dat_o[21] = net168;
 assign wbs_dat_o[22] = net169;
 assign wbs_dat_o[23] = net170;
 assign wbs_dat_o[24] = net171;
 assign wbs_dat_o[25] = net172;
 assign wbs_dat_o[26] = net173;
 assign wbs_dat_o[27] = net174;
 assign wbs_dat_o[28] = net175;
 assign wbs_dat_o[29] = net176;
 assign wbs_dat_o[2] = net149;
 assign wbs_dat_o[30] = net177;
 assign wbs_dat_o[31] = net178;
 assign wbs_dat_o[3] = net150;
 assign wbs_dat_o[4] = net151;
 assign wbs_dat_o[5] = net152;
 assign wbs_dat_o[6] = net153;
 assign wbs_dat_o[7] = net154;
 assign wbs_dat_o[8] = net155;
 assign wbs_dat_o[9] = net156;
endmodule

