* NGSPICE file created from tiny_user_project.ext - technology: gf180mcuC

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fill_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fill_2 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_4 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fill_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fill_1 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__antenna abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__antenna I VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dffq_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dffq_1 D CLK Q VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__mux2_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__mux2_2 I0 I1 S Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__buf_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__buf_1 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_8 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_8 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai21_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai21_1 A1 A2 B ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor2_1 A1 A2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_64 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_64 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__filltie abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__filltie VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_32 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_32 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand2_1 A1 A2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi21_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi21_1 A1 A2 B ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi22_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi22_1 A1 A2 B1 B2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi21_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi21_2 A1 A2 B ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 D RN CLK Q VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__mux4_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__mux4_1 I0 I1 I2 I3 S0 S1 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__xnor2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__xnor2_1 A1 A2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand3_1 A1 A2 A3 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_16 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_16 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai22_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai22_1 A1 A2 B1 B2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkinv_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkinv_1 I ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__buf_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__buf_2 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand2_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand2_2 A1 A2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__tiel abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__tiel ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai211_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai211_1 A1 A2 B C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand3_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand3_2 A1 A2 A3 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai221_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai221_1 A1 A2 B1 B2 C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__and3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__and3_1 A1 A2 A3 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__xor2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__xor2_1 A1 A2 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkinv_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkinv_2 I ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__endcap abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__endcap VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__xor3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__xor3_1 A1 A2 A3 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__and2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__and2_1 A1 A2 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi221_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi221_1 A1 A2 B1 B2 C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand3_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand3_4 A1 A2 A3 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi222_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi222_1 A1 A2 B1 B2 C1 C2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__or3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__or3_1 A1 A2 A3 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai211_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai211_4 A1 A2 B C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__inv_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__inv_1 I ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__and4_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__and4_1 A1 A2 A3 A4 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai31_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai31_1 A1 A2 A3 B ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi22_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi22_2 A1 A2 B1 B2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai211_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai211_2 A1 A2 B C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand4_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand4_1 A1 A2 A3 A4 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor3_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor3_2 A1 A2 A3 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi221_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi221_2 A1 A2 B1 B2 C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi211_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi211_2 A1 A2 B C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor3_1 A1 A2 A3 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__or2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__or2_1 A1 A2 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi211_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi211_1 A1 A2 B C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai32_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai32_1 A1 A2 A3 B1 B2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__tieh abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__tieh Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai21_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai21_2 A1 A2 B ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai221_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai221_2 A1 A2 B1 B2 C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor4_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor4_1 A1 A2 A3 A4 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand4_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand4_2 A1 A2 A3 A4 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__xnor3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__xnor3_1 A1 A2 A3 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor4_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor4_4 A1 A2 A3 A4 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__buf_20 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__buf_20 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai222_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai222_1 A1 A2 B1 B2 C1 C2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi221_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi221_4 A1 A2 B1 B2 C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi211_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi211_4 A1 A2 B C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor4_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor4_2 A1 A2 A3 A4 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor2_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor2_2 A1 A2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai222_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai222_4 A1 A2 B1 B2 C1 C2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai22_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai22_2 A1 A2 B1 B2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai32_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai32_2 A1 A2 A3 B1 B2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi22_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi22_4 A1 A2 B1 B2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dffrnq_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dffrnq_2 D RN CLK Q VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai33_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai33_1 A1 A2 A3 B1 B2 B3 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai221_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai221_4 A1 A2 B1 B2 C ZN VDD VSS
.ends

.subckt tiny_user_project io_in[0] io_in[10] io_in[11] io_in[12] io_in[13] io_in[14]
+ io_in[15] io_in[16] io_in[17] io_in[18] io_in[19] io_in[1] io_in[20] io_in[21] io_in[22]
+ io_in[23] io_in[24] io_in[25] io_in[26] io_in[27] io_in[28] io_in[29] io_in[2] io_in[30]
+ io_in[31] io_in[32] io_in[33] io_in[34] io_in[35] io_in[36] io_in[37] io_in[3] io_in[4]
+ io_in[5] io_in[6] io_in[7] io_in[8] io_in[9] io_oeb[0] io_oeb[10] io_oeb[11] io_oeb[12]
+ io_oeb[13] io_oeb[14] io_oeb[15] io_oeb[16] io_oeb[17] io_oeb[18] io_oeb[19] io_oeb[1]
+ io_oeb[20] io_oeb[21] io_oeb[22] io_oeb[23] io_oeb[24] io_oeb[25] io_oeb[26] io_oeb[27]
+ io_oeb[28] io_oeb[29] io_oeb[2] io_oeb[30] io_oeb[31] io_oeb[32] io_oeb[33] io_oeb[34]
+ io_oeb[35] io_oeb[36] io_oeb[37] io_oeb[3] io_oeb[4] io_oeb[5] io_oeb[6] io_oeb[7]
+ io_oeb[8] io_oeb[9] io_out[0] io_out[10] io_out[11] io_out[12] io_out[13] io_out[14]
+ io_out[15] io_out[16] io_out[17] io_out[18] io_out[19] io_out[1] io_out[20] io_out[21]
+ io_out[22] io_out[23] io_out[24] io_out[25] io_out[26] io_out[27] io_out[28] io_out[29]
+ io_out[2] io_out[30] io_out[31] io_out[32] io_out[33] io_out[34] io_out[35] io_out[36]
+ io_out[37] io_out[3] io_out[4] io_out[5] io_out[6] io_out[7] io_out[8] io_out[9]
+ la_data_in[0] la_data_in[10] la_data_in[11] la_data_in[12] la_data_in[13] la_data_in[14]
+ la_data_in[15] la_data_in[16] la_data_in[17] la_data_in[18] la_data_in[19] la_data_in[1]
+ la_data_in[20] la_data_in[21] la_data_in[22] la_data_in[23] la_data_in[24] la_data_in[25]
+ la_data_in[26] la_data_in[27] la_data_in[28] la_data_in[29] la_data_in[2] la_data_in[30]
+ la_data_in[31] la_data_in[32] la_data_in[33] la_data_in[34] la_data_in[35] la_data_in[36]
+ la_data_in[37] la_data_in[38] la_data_in[39] la_data_in[3] la_data_in[40] la_data_in[41]
+ la_data_in[42] la_data_in[43] la_data_in[44] la_data_in[45] la_data_in[46] la_data_in[47]
+ la_data_in[48] la_data_in[49] la_data_in[4] la_data_in[50] la_data_in[51] la_data_in[52]
+ la_data_in[53] la_data_in[54] la_data_in[55] la_data_in[56] la_data_in[57] la_data_in[58]
+ la_data_in[59] la_data_in[5] la_data_in[60] la_data_in[61] la_data_in[62] la_data_in[63]
+ la_data_in[6] la_data_in[7] la_data_in[8] la_data_in[9] la_data_out[0] la_data_out[10]
+ la_data_out[11] la_data_out[12] la_data_out[13] la_data_out[14] la_data_out[15]
+ la_data_out[16] la_data_out[17] la_data_out[18] la_data_out[19] la_data_out[1] la_data_out[20]
+ la_data_out[21] la_data_out[22] la_data_out[23] la_data_out[24] la_data_out[25]
+ la_data_out[26] la_data_out[27] la_data_out[28] la_data_out[29] la_data_out[2] la_data_out[30]
+ la_data_out[31] la_data_out[32] la_data_out[33] la_data_out[34] la_data_out[35]
+ la_data_out[36] la_data_out[37] la_data_out[38] la_data_out[39] la_data_out[3] la_data_out[40]
+ la_data_out[41] la_data_out[42] la_data_out[43] la_data_out[44] la_data_out[45]
+ la_data_out[46] la_data_out[47] la_data_out[48] la_data_out[49] la_data_out[4] la_data_out[50]
+ la_data_out[51] la_data_out[52] la_data_out[53] la_data_out[54] la_data_out[55]
+ la_data_out[56] la_data_out[57] la_data_out[58] la_data_out[59] la_data_out[5] la_data_out[60]
+ la_data_out[61] la_data_out[62] la_data_out[63] la_data_out[6] la_data_out[7] la_data_out[8]
+ la_data_out[9] la_oenb[0] la_oenb[10] la_oenb[11] la_oenb[12] la_oenb[13] la_oenb[14]
+ la_oenb[15] la_oenb[16] la_oenb[17] la_oenb[18] la_oenb[19] la_oenb[1] la_oenb[20]
+ la_oenb[21] la_oenb[22] la_oenb[23] la_oenb[24] la_oenb[25] la_oenb[26] la_oenb[27]
+ la_oenb[28] la_oenb[29] la_oenb[2] la_oenb[30] la_oenb[31] la_oenb[32] la_oenb[33]
+ la_oenb[34] la_oenb[35] la_oenb[36] la_oenb[37] la_oenb[38] la_oenb[39] la_oenb[3]
+ la_oenb[40] la_oenb[41] la_oenb[42] la_oenb[43] la_oenb[44] la_oenb[45] la_oenb[46]
+ la_oenb[47] la_oenb[48] la_oenb[49] la_oenb[4] la_oenb[50] la_oenb[51] la_oenb[52]
+ la_oenb[53] la_oenb[54] la_oenb[55] la_oenb[56] la_oenb[57] la_oenb[58] la_oenb[59]
+ la_oenb[5] la_oenb[60] la_oenb[61] la_oenb[62] la_oenb[63] la_oenb[6] la_oenb[7]
+ la_oenb[8] la_oenb[9] user_clock2 user_irq[0] user_irq[1] user_irq[2] vdd vss wb_clk_i
+ wb_rst_i wbs_ack_o wbs_adr_i[0] wbs_adr_i[10] wbs_adr_i[11] wbs_adr_i[12] wbs_adr_i[13]
+ wbs_adr_i[14] wbs_adr_i[15] wbs_adr_i[16] wbs_adr_i[17] wbs_adr_i[18] wbs_adr_i[19]
+ wbs_adr_i[1] wbs_adr_i[20] wbs_adr_i[21] wbs_adr_i[22] wbs_adr_i[23] wbs_adr_i[24]
+ wbs_adr_i[25] wbs_adr_i[26] wbs_adr_i[27] wbs_adr_i[28] wbs_adr_i[29] wbs_adr_i[2]
+ wbs_adr_i[30] wbs_adr_i[31] wbs_adr_i[3] wbs_adr_i[4] wbs_adr_i[5] wbs_adr_i[6]
+ wbs_adr_i[7] wbs_adr_i[8] wbs_adr_i[9] wbs_cyc_i wbs_dat_i[0] wbs_dat_i[10] wbs_dat_i[11]
+ wbs_dat_i[12] wbs_dat_i[13] wbs_dat_i[14] wbs_dat_i[15] wbs_dat_i[16] wbs_dat_i[17]
+ wbs_dat_i[18] wbs_dat_i[19] wbs_dat_i[1] wbs_dat_i[20] wbs_dat_i[21] wbs_dat_i[22]
+ wbs_dat_i[23] wbs_dat_i[24] wbs_dat_i[25] wbs_dat_i[26] wbs_dat_i[27] wbs_dat_i[28]
+ wbs_dat_i[29] wbs_dat_i[2] wbs_dat_i[30] wbs_dat_i[31] wbs_dat_i[3] wbs_dat_i[4]
+ wbs_dat_i[5] wbs_dat_i[6] wbs_dat_i[7] wbs_dat_i[8] wbs_dat_i[9] wbs_dat_o[0] wbs_dat_o[10]
+ wbs_dat_o[11] wbs_dat_o[12] wbs_dat_o[13] wbs_dat_o[14] wbs_dat_o[15] wbs_dat_o[16]
+ wbs_dat_o[17] wbs_dat_o[18] wbs_dat_o[19] wbs_dat_o[1] wbs_dat_o[20] wbs_dat_o[21]
+ wbs_dat_o[22] wbs_dat_o[23] wbs_dat_o[24] wbs_dat_o[25] wbs_dat_o[26] wbs_dat_o[27]
+ wbs_dat_o[28] wbs_dat_o[29] wbs_dat_o[2] wbs_dat_o[30] wbs_dat_o[31] wbs_dat_o[3]
+ wbs_dat_o[4] wbs_dat_o[5] wbs_dat_o[6] wbs_dat_o[7] wbs_dat_o[8] wbs_dat_o[9] wbs_sel_i[0]
+ wbs_sel_i[1] wbs_sel_i[2] wbs_sel_i[3] wbs_stb_i wbs_we_i
XFILLER_39_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8507__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6209__A2 _1781_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7257__I1 _3312_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_726 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_748 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7963_ _0189_ net1 mod.Data_Mem.F_M.MRAM\[779\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_82_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7009__I1 mod.Data_Mem.F_M.MRAM\[17\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6914_ _3253_ mod.Data_Mem.F_M.MRAM\[13\]\[5\] _3381_ _3383_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_78_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7894_ _0120_ net1 mod.Data_Mem.F_M.MRAM\[27\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_165_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_1194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6845_ _3256_ mod.Data_Mem.F_M.MRAM\[769\]\[6\] _3340_ _3345_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_74_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_168_29 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6776_ _3297_ _3298_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_23_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5196__A2 _1825_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3988_ _0664_ _0665_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_50_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_8515_ _0019_ net1 mod.Data_Mem.F_M.out_data\[59\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__8499__D _0003_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5727_ _2209_ _2352_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__7256__I _3584_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_148_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8446_ _0542_ net1 mod.Data_Mem.F_M.MRAM\[793\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5658_ _2288_ mod.Data_Mem.F_M.MRAM\[796\]\[2\] _2268_ _2289_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_50_1080 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4609_ _1201_ _1257_ _1280_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_164_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_8377_ _0473_ net1 mod.Data_Mem.F_M.MRAM\[784\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_102_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5743__I1 mod.Data_Mem.F_M.MRAM\[3\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5589_ _1549_ _2226_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__8037__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_117_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7328_ _3297_ _3634_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5932__C _2552_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_753 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8126__RN net2 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6448__A2 _3054_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7259_ mod.Data_Mem.F_M.MRAM\[31\]\[5\] _3316_ _3590_ _3592_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_85_1198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4459__A1 _1125_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_133_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8187__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7248__I1 _3293_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3202 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3213 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_895 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3224 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3235 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2501 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3246 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3257 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2512 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3959__I _0635_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2523 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2534 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2545 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1800 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_165_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2556 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1811 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1822 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2567 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_781 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2578 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1833 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2589 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_943 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1844 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1855 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3985__A3 mod.Arithmetic.CN.I_in\[64\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1866 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_158_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_42_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1877 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1888 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6384__A1 _2134_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5187__A2 mod.Data_Mem.F_M.MRAM\[771\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1899 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6384__B2 _2216_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5982__I1 mod.Data_Mem.F_M.MRAM\[771\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6070__I _2686_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_761 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5734__I1 mod.Data_Mem.F_M.MRAM\[15\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4698__A1 _0620_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_1216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8117__RN net2 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7487__I1 mod.Data_Mem.F_M.MRAM\[781\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5414__I _1725_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_615 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_81 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_748 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_91_320 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6998__I0 _3395_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4960_ _1625_ _1628_ _1629_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_33_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4891_ _1547_ _1552_ _1559_ _1560_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_71_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6630_ _3205_ _0106_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6375__A1 _2779_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_784 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_80_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_6561_ mod.Data_Mem.F_M.MRAM\[781\]\[7\] _2596_ _3023_ mod.Data_Mem.F_M.MRAM\[769\]\[7\]
+ _3163_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_164_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_8300_ _0396_ net1 mod.Data_Mem.F_M.MRAM\[773\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5512_ _2151_ mod.Data_Mem.F_M.MRAM\[30\]\[7\] _2153_ _2154_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XANTENNA__6127__A1 _1726_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_536 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6492_ _2511_ mod.Data_Mem.F_M.MRAM\[0\]\[4\] _2103_ _3097_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_69_1116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_8231_ mod.P1.instr_reg\[17\] net2 net1 mod.P2.dest_reg1\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_69_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5443_ _1548_ _2092_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_146_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_133_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_160_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8162_ mod.Data_Mem.F_M.out_data\[72\] net2 net1 mod.Arithmetic.I_out\[72\] vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_5374_ _2032_ _2033_ _2034_ _2035_ _1844_ _1642_ _2036_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__4153__A3 mod.Arithmetic.CN.I_in\[33\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7113_ _3504_ _0290_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__7478__I1 mod.Data_Mem.F_M.MRAM\[780\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8108__RN net2 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4325_ _0994_ _0998_ _0999_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_8093_ mod.Data_Mem.F_M.out_data\[3\] net2 net1 mod.Arithmetic.ACTI.x\[3\] vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_99_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7044_ _3468_ _0257_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_87_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4256_ _0621_ _0930_ _0658_ _0931_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_68_840 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4187_ _0802_ _0818_ _0862_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_28_726 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6989__I0 _3405_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_1109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_17 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1107 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_7946_ _0172_ net1 mod.Data_Mem.F_M.MRAM\[789\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1129 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_7877_ _0103_ net1 mod.Data_Mem.F_M.MRAM\[24\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_51_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_464 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_773 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6828_ mod.Data_Mem.F_M.dest\[1\] _3333_ _3334_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__6366__A1 _1941_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_1180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6759_ _3286_ _0154_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_104_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_1153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6118__A1 _2373_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7166__I0 _3537_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_1216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5943__B _2563_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_163_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_152_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8429_ _0525_ net1 mod.Data_Mem.F_M.MRAM\[791\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_3_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_285 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_981 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3010 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3021 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3032 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3043 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_18_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3054 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2320 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6065__I _2681_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3065 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3076 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2331 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3087 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2342 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3098 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2353 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2364 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2375 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1630 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1641 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_148_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2386 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2397 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1652 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_159_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1674 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6357__A1 _2904_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8202__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1685 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_784 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1696 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_105_1007 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_1018 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_169_72 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_30_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4907__A2 _1575_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_146_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_127_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6109__A1 _2692_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7157__I0 _3531_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5580__A2 mod.Data_Mem.F_M.MRAM\[30\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8352__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_539 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_1002 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4110_ _0781_ _0780_ _0785_ _0786_ _0787_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_69_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5090_ _1756_ _1757_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_69_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6293__B1 mod.Data_Mem.F_M.MRAM\[14\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4983__I _1561_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4041_ mod.Arithmetic.I_out\[72\] _0718_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__5080__S _1746_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_640 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7800_ _3898_ _0583_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_92_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5992_ _2560_ _2611_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_64_397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7731_ _3859_ _0553_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4943_ _1567_ _1612_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_127_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6703__I net8 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5747__C _1498_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7662_ mod.Data_Mem.F_M.MRAM\[790\]\[7\] _3825_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4874_ _1542_ _1543_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_20_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_1197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6613_ mod.Data_Mem.F_M.MRAM\[24\]\[2\] _3197_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_7593_ _3786_ _3787_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__5020__A1 _1686_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_165_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_20_467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6544_ _3145_ _3146_ _2474_ _3147_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__7148__I0 _3523_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_145_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_355 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6475_ _3004_ _3080_ _3081_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_134_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5859__B1 _2478_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8214_ _0315_ net1 mod.Data_Mem.F_M.MRAM\[22\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_161_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5426_ _2067_ _2082_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6520__A1 _3106_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5323__A2 _1673_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6371__I1 _2035_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8145_ mod.Data_Mem.F_M.out_data\[55\] net2 net1 mod.Arithmetic.CN.I_in\[55\] vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_5357_ mod.Data_Mem.F_M.MRAM\[799\]\[6\] _1913_ _2019_ _2020_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__7470__S _3707_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4308_ _0980_ _0981_ _0982_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_88_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8076_ mod.P3.Res\[4\] net2 net1 net7 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XANTENNA__7320__I0 _3615_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5288_ mod.Data_Mem.F_M.MRAM\[775\]\[5\] mod.Data_Mem.F_M.MRAM\[774\]\[5\] _1951_
+ _1952_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__4893__I _1561_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7027_ _3447_ _3457_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_4239_ _0615_ mod.Arithmetic.CN.I_in\[66\] _0914_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_68_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6036__B1 _2536_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5003__B _1668_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8225__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_167_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_55_397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7929_ _0155_ net1 mod.Data_Mem.F_M.MRAM\[8\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_43_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_356 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6339__A1 _2779_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8375__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5011__A1 _1677_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4133__I _0808_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7139__I0 _3508_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_1051 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5392__C _1822_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6511__A1 _2587_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_151_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_140_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_105_561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_78_467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_78_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_898 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_1017 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_1148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2150 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5848__B _2429_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2161 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2172 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2183 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2194 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1460 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1471 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1482 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_8518__184 net184 vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_9_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_147_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4590_ _1260_ _1261_ _1262_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_70_1072 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5553__A2 _2185_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_31_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_6_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6260_ _2706_ _2873_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_6_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5211_ mod.Data_Mem.F_M.MRAM\[7\]\[4\] mod.Data_Mem.F_M.MRAM\[6\]\[4\] _1875_ _1876_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_43_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7892__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6191_ _1661_ _2804_ _2805_ _2763_ _2806_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_69_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5142_ mod.Data_Mem.F_M.MRAM\[5\]\[3\] mod.Data_Mem.F_M.MRAM\[4\]\[3\] _1510_ _1808_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_97_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5069__A1 _1734_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5073_ _1738_ _1739_ _1562_ _1740_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_84_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8248__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5864__I0 mod.Data_Mem.F_M.MRAM\[18\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4024_ _0696_ mod.Arithmetic.I_out\[78\] _0697_ _0701_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_84_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4292__A2 _0878_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4218__I mod.Arithmetic.CN.I_in\[34\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6569__A1 _0612_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8398__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5975_ _2531_ _2586_ _2594_ _2595_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_80_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4662__B _1251_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7714_ mod.Data_Mem.F_M.MRAM\[794\]\[1\] _3851_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4926_ _1492_ _1595_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_33_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7645_ _3816_ _0510_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4857_ _1525_ _1526_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_14_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7576_ _3749_ mod.Data_Mem.F_M.MRAM\[785\]\[2\] _3773_ _3776_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4788_ _1234_ _1344_ _1458_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_101_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6527_ _3111_ _3130_ _3131_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_119_675 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_84_1208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6458_ _2063_ _3064_ _3065_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_122_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_133_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4355__I0 _0775_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5409_ _2063_ _0010_ _0008_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_121_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6389_ mod.Data_Mem.F_M.MRAM\[781\]\[7\] _2901_ _2902_ mod.Data_Mem.F_M.MRAM\[780\]\[7\]
+ _2998_ _2999_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_88_710 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_1000 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_8128_ mod.Data_Mem.F_M.out_data\[38\] net2 net1 mod.Arithmetic.CN.I_in\[38\] vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_47_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8059_ _0268_ net1 mod.Data_Mem.F_M.MRAM\[20\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_87_264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_56_651 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5480__A1 _1803_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4128__I _0803_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_879 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4586__A3 _1257_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5783__A2 _2407_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_169_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_1056 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6032__I0 mod.Data_Mem.F_M.MRAM\[784\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_169_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_156_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7780__I0 _3784_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_109_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5299__A1 _1631_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_1016 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_1185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_765 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_94_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_152_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_895 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5422__I _2079_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_19_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8540__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4038__I mod.Arithmetic.CN.I_in\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_610 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_37_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7763__A3 _3371_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6253__I _2374_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5760_ _1840_ _2385_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_15_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5774__A2 mod.Data_Mem.F_M.MRAM\[789\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4711_ _1369_ _1381_ _1382_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XTAP_1290 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5691_ _2319_ mod.Data_Mem.F_M.MRAM\[797\]\[4\] _2320_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__7285__S _3606_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7430_ _3688_ _0423_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4642_ _1063_ _1178_ mod.Arithmetic.CN.I_in\[30\] _1313_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_30_584 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7361_ mod.Data_Mem.F_M.MRAM\[772\]\[5\] _3654_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4573_ _1125_ _1244_ _1245_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_116_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6312_ _2870_ _1950_ _2924_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_7292_ _3305_ _3612_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5129__I2 _1789_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_104_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6243_ _2853_ _2856_ _2743_ _2857_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_131_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8070__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5385__S1 _2009_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_6174_ _1898_ _2789_ _2790_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_130_158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_85_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5125_ mod.Data_Mem.F_M.MRAM\[784\]\[2\] _1792_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_97_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_131_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5056_ mod.Data_Mem.F_M.src\[8\] _1724_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_73_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5462__A1 _2108_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2908 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4007_ mod.Arithmetic.CN.I_in\[17\] _0684_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_84_278 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2919 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_429 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_25_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_643 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_168_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_129_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5958_ mod.Data_Mem.F_M.MRAM\[18\]\[5\] mod.Data_Mem.F_M.MRAM\[19\]\[5\] _2161_ _2578_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_80_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_52_197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4909_ _1502_ _1578_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_5889_ _1707_ _2511_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_166_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_7628_ _3319_ _3798_ _3808_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_138_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_461 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6190__A2 _1731_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7559_ _3765_ mod.Data_Mem.F_M.MRAM\[784\]\[3\] _3760_ _3766_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_14_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8413__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_1152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_162_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_1196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_161_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_150_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_122_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8563__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4256__A2 _0930_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_749 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_28_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_147_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_974 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_44_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_1009 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5508__A2 _2148_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_157_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_23 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_32_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5417__I _2075_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6181__A2 _2795_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8093__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4192__A1 _0623_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7505__I0 _3731_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_113_615 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7632__I mod.Data_Mem.F_M.MRAM\[788\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5353__S _1580_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5367__S1 _1590_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5141__B1 _1730_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_348 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_359 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4495__A2 _1072_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_584 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7930__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5444__A1 _2092_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5295__I1 _1952_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_278 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6930_ _3394_ _0217_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_35_610 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5995__A2 mod.Data_Mem.F_M.MRAM\[786\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_930 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6861_ mod.Data_Mem.F_M.MRAM\[779\]\[6\] _3353_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__7197__A1 _3555_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_985 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6912__S _3381_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5812_ _2152_ mod.Data_Mem.F_M.MRAM\[771\]\[1\] _2436_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6792_ _3310_ _0163_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_34_197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5743_ mod.Data_Mem.F_M.MRAM\[2\]\[0\] mod.Data_Mem.F_M.MRAM\[3\]\[0\] _1515_ _2368_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_8531_ _0035_ net1 mod.Data_Mem.F_M.out_data\[43\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_148_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6711__I net10 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8436__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8462_ _0558_ net1 mod.Data_Mem.F_M.MRAM\[795\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5674_ _2300_ _2303_ _2304_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_30_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7413_ mod.Data_Mem.F_M.MRAM\[775\]\[7\] _3680_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4625_ _1292_ _1295_ _1296_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_8393_ _0489_ net1 mod.Data_Mem.F_M.MRAM\[786\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__6172__A2 _1684_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7344_ _3315_ _3645_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_144_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4556_ _0645_ mod.Arithmetic.CN.I_in\[53\] _1114_ _1116_ _1228_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__8586__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7275_ mod.Data_Mem.F_M.MRAM\[5\]\[5\] _3600_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4487_ _1089_ _1102_ _1159_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_143_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_968 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6226_ _1585_ _2839_ _2840_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_44_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_1082 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6157_ _2425_ mod.Data_Mem.F_M.MRAM\[22\]\[1\] mod.Data_Mem.F_M.MRAM\[23\]\[1\] _2188_
+ _2773_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_860 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_724 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_1093 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_871 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5062__I _1537_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_893 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5108_ _1598_ _1775_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_85_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6088_ _2012_ _1610_ _2705_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_100_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5435__A1 _2063_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2705 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5039_ _1567_ _1707_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_122_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2716 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_66_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2727 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2738 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2749 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_90_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_167_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_51_1037 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4961__A3 _1560_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_110_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__4174__A1 _0825_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_108_987 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_108_998 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput7 net7 io_out[20] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XFILLER_134_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7953__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_1111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4477__A2 _0716_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5901__S _2522_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_746 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_1188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8309__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_749 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5977__A2 mod.Data_Mem.F_M.MRAM\[783\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_974 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_985 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_782 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8459__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5729__A2 _1553_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_160_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_170 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_181 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_118_718 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6154__A2 _1659_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5147__I _1517_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7563__S _3760_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4410_ _1048_ _1077_ _1082_ _1083_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
X_5390_ mod.Data_Mem.F_M.MRAM\[785\]\[7\] mod.Data_Mem.F_M.MRAM\[784\]\[7\] _1813_
+ _2052_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_126_751 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4704__A3 _1125_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_1022 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4341_ _1008_ _1014_ _1015_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_153_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_125_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_98_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7060_ mod.Data_Mem.F_M.MRAM\[20\]\[1\] _3477_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_114_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4272_ _0867_ _0885_ _0946_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_67_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_819 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6701__I1 mod.Data_Mem.F_M.MRAM\[28\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_1211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6011_ _2379_ _2618_ _2625_ _2626_ _2629_ _2630_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XANTENNA__5665__A1 _2295_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4468__A2 _1108_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6907__S _3376_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7962_ _0188_ net1 mod.Data_Mem.F_M.MRAM\[779\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6913_ _3382_ _0212_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_7893_ _0119_ net1 mod.Data_Mem.F_M.MRAM\[25\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_51_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_911 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4640__A2 _0679_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_1015 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6844_ _1955_ _3337_ _3344_ _0181_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_23_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_432 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4670__B _1340_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6775_ mod.Data_Mem.F_M.dest\[8\] mod.DMen_reg2 _3297_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__6393__A2 _3002_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5196__A3 _1861_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3987_ _0633_ mod.Arithmetic.ACTI.x\[0\] _0664_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__8071__RN net2 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6441__I _2092_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_149_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_8514_ _0018_ net1 mod.Data_Mem.F_M.out_data\[58\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5726_ _2351_ _0055_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__5028__S0 _1695_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_718 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8445_ _0541_ net1 mod.Data_Mem.F_M.MRAM\[793\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5657_ _1609_ _2288_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__5057__I _1724_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7473__S _3707_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4156__A1 _0657_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7976__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_1092 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4608_ _1159_ _1196_ _1278_ _1279_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_117_751 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8376_ _0472_ net1 mod.Data_Mem.F_M.MRAM\[784\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5588_ _1800_ _2158_ _2093_ _2225_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_117_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4896__I _1564_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7327_ _3633_ _0375_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_2_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4539_ _1209_ _1210_ _1211_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_137_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_1155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7258_ _3591_ _0348_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_120_916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_77_307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5656__A1 _2151_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6209_ _2186_ _1781_ _2824_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_131_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7189_ _3523_ mod.Data_Mem.F_M.MRAM\[29\]\[0\] _3550_ _3551_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_58_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_852 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_690 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3203 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_133_55 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_3214 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3225 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3236 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3247 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2502 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5520__I _1942_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5959__A2 _2578_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3258 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2513 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2524 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2535 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2546 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1801 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2557 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1812 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2568 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1823 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2579 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1834 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_1845 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1856 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1867 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1878 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1889 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_988 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6384__A2 mod.Data_Mem.F_M.MRAM\[15\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5395__C _1629_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_690 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_166_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_154_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_5_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_927 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5647__A1 _2168_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8131__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_151_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_68_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_690 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5430__I _2084_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6998__I1 mod.Data_Mem.F_M.MRAM\[17\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8281__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_149_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_64_568 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4890_ mod.Data_Mem.F_M.MRAM\[15\]\[0\] _1536_ mod.Data_Mem.F_M.MRAM\[31\]\[0\] _1558_
+ _1551_ _1559_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_20_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_796 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4386__A1 _0806_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7999__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6560_ _2831_ _3161_ _3162_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_158_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5511_ _2152_ mod.Data_Mem.F_M.MRAM\[31\]\[7\] _2153_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_73_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6491_ _2728_ mod.Data_Mem.F_M.MRAM\[1\]\[4\] _3096_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_160_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4138__A1 _0813_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8230_ mod.P1.instr_reg\[13\] net2 net1 mod.P2.dest_reg1\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_5442_ _2008_ _2091_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_69_1128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4689__A2 _1354_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5373_ mod.Data_Mem.F_M.MRAM\[17\]\[7\] mod.Data_Mem.F_M.MRAM\[16\]\[7\] _1894_ _2035_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_8161_ mod.Data_Mem.F_M.out_data\[71\] net2 net1 mod.Arithmetic.CN.I_in\[71\] vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XANTENNA__6210__B _2739_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7112_ _3452_ mod.Data_Mem.F_M.MRAM\[3\]\[2\] _3501_ _3504_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4324_ _0930_ _0995_ _0996_ _0997_ _0998_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
X_8092_ mod.Data_Mem.F_M.out_data\[2\] net2 net1 mod.Arithmetic.ACTI.x\[2\] vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XANTENNA__5638__A1 _2270_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7043_ _3450_ mod.Data_Mem.F_M.MRAM\[1\]\[1\] _3466_ _3468_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_113_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4255_ mod.Arithmetic.CN.I_in\[49\] _0930_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_87_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_949 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4186_ _0801_ _0852_ _0861_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_80_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_682 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_27_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_535 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6989__I1 mod.Data_Mem.F_M.MRAM\[16\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6063__A1 _2534_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6063__B2 _2414_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7945_ _0171_ net1 mod.Data_Mem.F_M.MRAM\[789\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_36_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1108 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1119 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4613__A2 _1187_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7468__S _3707_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_169_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7876_ _0102_ net1 mod.Data_Mem.F_M.MRAM\[24\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6827_ mod.Data_Mem.F_M.dest\[0\] _3333_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__8004__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_1121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_137_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6758_ mod.Data_Mem.F_M.MRAM\[8\]\[2\] _3286_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_91_1192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_109_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5709_ _2315_ mod.Data_Mem.F_M.MRAM\[28\]\[6\] _2316_ _2336_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_148_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6118__A2 _2687_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7166__I1 mod.Data_Mem.F_M.MRAM\[12\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6689_ _3241_ _0129_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_87_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8428_ _0524_ net1 mod.Data_Mem.F_M.MRAM\[791\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_164_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_124_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8154__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_77 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_88 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_8359_ _0455_ net1 mod.Data_Mem.F_M.MRAM\[781\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_2_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_105_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_160_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_24_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4301__A1 _0901_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3000 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_59_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_822 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3011 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3022 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3033 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3044 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3055 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2310 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_34_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3066 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2321 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3077 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2332 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2343 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3088 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_1010 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4604__A2 _1258_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3099 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2354 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2365 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1620 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2376 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_730 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1631 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2387 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1642 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2398 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1653 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1664 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1675 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7177__I mod.Data_Mem.F_M.MRAM\[22\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6357__A2 mod.Data_Mem.F_M.MRAM\[783\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__7554__A1 _3610_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1686 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6081__I _1756_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1697 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4368__A1 _0901_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5565__B1 mod.Data_Mem.F_M.MRAM\[31\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_168_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_167_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_1161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4540__A1 _1208_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_155_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_1069 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7640__I mod.Data_Mem.F_M.MRAM\[788\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_150_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_111_757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6293__A1 _2904_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4040_ _0710_ _0712_ _0714_ _0716_ _0717_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__5340__I0 mod.Data_Mem.F_M.MRAM\[771\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_822 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6256__I _2686_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5160__I _1663_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5991_ _2414_ _2595_ _2610_ _0061_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_80_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7730_ mod.Data_Mem.F_M.MRAM\[795\]\[1\] _3859_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__8027__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_1132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4942_ _1608_ _1610_ _1611_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_162_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_33_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7661_ _3824_ _0518_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_21_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4873_ _1541_ _1542_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6612_ _3196_ _0097_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4359__A1 _0781_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7592_ _3604_ _3446_ _3758_ _3786_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_4
XANTENNA__8177__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_159_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6543_ _3106_ mod.Data_Mem.F_M.MRAM\[769\]\[6\] _3107_ _3146_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__7148__I1 mod.Data_Mem.F_M.MRAM\[12\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6474_ _3026_ _2304_ _3006_ _2523_ _2529_ _2510_ _3080_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_146_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_106_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5859__A1 _2435_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8213_ _0314_ net1 mod.Data_Mem.F_M.MRAM\[22\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_106_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_160_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5425_ _2081_ _0010_ _0016_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__6520__A2 mod.Data_Mem.F_M.MRAM\[781\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5356_ _2011_ _2018_ _1775_ _2019_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_99_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8144_ mod.Data_Mem.F_M.out_data\[54\] net2 net1 mod.Arithmetic.CN.I_in\[54\] vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_114_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4307_ _0893_ _0829_ _0892_ mod.Arithmetic.CN.I_in\[33\] _0981_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
X_8075_ mod.P3.Res\[3\] net2 net1 net6 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_87_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5287_ _1816_ _1951_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_101_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7550__I _3759_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7026_ _3248_ _3456_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4238_ _0842_ _0911_ _0912_ _0913_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or3_1
XFILLER_56_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_822 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5070__I _1606_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4169_ _0844_ mod.Arithmetic.ACTI.x\[1\] _0845_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_83_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6036__B2 _2649_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5003__C _1670_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_83_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_23 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7928_ _0154_ net1 mod.Data_Mem.F_M.MRAM\[8\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_93_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_169_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_169_713 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_54_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_70_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7859_ _3913_ _3917_ _0608_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_11_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5954__B _2075_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4070__I0 _0630_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_149_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7139__I1 mod.Data_Mem.F_M.MRAM\[19\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5673__C _2268_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4770__A1 _0624_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_152_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_109_367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_165_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_136_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6511__A2 mod.Data_Mem.F_M.MRAM\[13\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_860 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_132_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6275__A1 _2872_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_63_1080 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_1121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6027__A1 _2416_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_1165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_73_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2140 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2151 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2162 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2173 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2184 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2195 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_159_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1461 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1472 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1483 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1494 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__4761__A1 _1285_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_115_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5210_ _1646_ _1875_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_6190_ _2761_ _1731_ _2805_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_130_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5141_ mod.Data_Mem.F_M.MRAM\[22\]\[3\] _1601_ _1730_ _1806_ _1507_ _1807_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_36_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_111_532 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5069__A2 _1735_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6266__A1 _2869_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5072_ mod.Data_Mem.F_M.MRAM\[3\]\[2\] mod.Data_Mem.F_M.MRAM\[2\]\[2\] _1647_ _1739_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_85_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_427 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5864__I1 mod.Data_Mem.F_M.MRAM\[19\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4023_ _0696_ mod.Arithmetic.I_out\[78\] _0697_ _0699_ _0700_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_4
XFILLER_84_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_855 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_65_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_1216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_983 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6569__A2 _3169_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_611 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5974_ _2410_ _2590_ _2593_ _2594_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_7713_ _3850_ _0544_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4925_ _1593_ _1594_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__7746__S _3867_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_7644_ mod.Data_Mem.F_M.MRAM\[788\]\[6\] _3816_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4856_ _1524_ _1525_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_20_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_165_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_7575_ _3775_ _0481_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4787_ _0624_ _1456_ _1457_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_20_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6526_ _2508_ _2333_ _3060_ _2605_ _2606_ _3107_ _3130_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_134_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_161_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6457_ mod.Data_Mem.F_M.MRAM\[13\]\[2\] _2382_ _2642_ mod.Data_Mem.F_M.MRAM\[1\]\[2\]
+ _3064_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_134_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4504__A1 _0806_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4355__I1 _0774_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5408_ _2068_ _0010_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6388_ _2903_ _2997_ _2998_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_121_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_893 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_138_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8127_ mod.Data_Mem.F_M.out_data\[37\] net2 net1 mod.Arithmetic.CN.I_in\[37\] vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_87_210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5339_ mod.Data_Mem.F_M.MRAM\[769\]\[6\] mod.Data_Mem.F_M.MRAM\[768\]\[6\] _1814_
+ _2002_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_87_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_852 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8058_ _0267_ net1 mod.Data_Mem.F_M.MRAM\[20\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_88_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7009_ _3405_ mod.Data_Mem.F_M.MRAM\[17\]\[7\] _3440_ _3444_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__5855__I1 mod.Data_Mem.F_M.MRAM\[783\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_169_1108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_28_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6009__A1 _2104_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5949__B _2568_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8342__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6804__I0 mod.Data_Mem.F_M.MRAM\[799\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_55_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5232__A2 _1896_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_1160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_169_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_571 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__4144__I mod.Arithmetic.CN.I_in\[32\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_157_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8492__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7780__I1 mod.Data_Mem.F_M.MRAM\[797\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4743__A1 mod.Arithmetic.CN.I_in\[47\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_153_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6496__A1 _2103_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_112_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_117_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5703__I _1581_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_83 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6248__A1 _2108_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_1197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_939 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_427 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7048__I0 _3454_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8229__RN net2 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_942 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_34_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6420__A1 _2184_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4054__I mod.Arithmetic.CN.I_in\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4710_ _1372_ _1380_ _1381_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_1291 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4982__A1 _1565_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5690_ _2096_ _2319_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_147_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6184__B1 mod.Data_Mem.F_M.MRAM\[15\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4641_ _1310_ _1311_ _1312_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_7360_ _3653_ _0388_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4572_ _0614_ mod.Arithmetic.ACTI.x\[5\] _1244_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_116_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_128_473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6311_ _2882_ _2921_ _2922_ _2884_ _2078_ _2923_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_143_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7291_ _1716_ _3609_ _3611_ _0361_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__5814__S _1918_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5129__I3 _1794_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8215__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6487__A1 _3004_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6242_ _2854_ _2855_ _2738_ _2856_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_89_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_1220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_157_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_131_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6173_ _2785_ _2786_ _2787_ _2788_ _2750_ _2789_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_69_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6239__A1 _2846_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5124_ _1790_ _1791_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_111_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8365__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5055_ mod.Data_Mem.F_M.MRAM\[783\]\[1\] _1699_ _1722_ _1723_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__5998__B1 _2616_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4006_ mod.Arithmetic.I_out\[74\] _0683_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XANTENNA__5462__A2 _2110_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2909 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_77_1002 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_1013 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_52_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_40_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5957_ _2534_ _2555_ _2577_ _2414_ _0060_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_52_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4908_ _1563_ _1570_ _1576_ _1577_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_33_390 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5888_ _2495_ _2510_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__7211__I0 _3527_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4899__I _1567_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7627_ _3807_ _0501_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4839_ _1507_ _1508_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__7275__I mod.Data_Mem.F_M.MRAM\[5\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7558_ _3308_ _3765_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_107_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6509_ _1491_ _3113_ _3114_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_88_1164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_1055 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_432 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7489_ _3638_ mod.Data_Mem.F_M.MRAM\[781\]\[1\] _3720_ _3722_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_49_1126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6478__A1 _2315_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_77 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_121_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_427 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5989__B1 _2602_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__3978__I _0654_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_1113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_17_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_71_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_71_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6402__A1 _2256_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7882__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_43_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_12_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_129_237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__8238__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6022__C _2091_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4192__A2 _0656_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7505__I1 mod.Data_Mem.F_M.MRAM\[781\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6469__A1 _2151_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_125_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8388__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5141__A1 mod.Data_Mem.F_M.MRAM\[22\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5141__B2 _1806_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_67_703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_1051 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_94_500 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4049__I _0691_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_950 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5295__I2 _1957_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_994 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6860_ _3352_ _0189_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_35_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_1208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7197__A2 _3550_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5811_ _2109_ _2435_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_34_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6791_ mod.Data_Mem.F_M.MRAM\[799\]\[3\] _3309_ _3300_ _3310_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_22_327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8530_ _0034_ net1 mod.Data_Mem.F_M.out_data\[42\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5742_ _2356_ _2367_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4955__A1 _1618_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_163_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8461_ _0557_ net1 mod.Data_Mem.F_M.MRAM\[795\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5673_ _2288_ mod.Data_Mem.F_M.MRAM\[28\]\[3\] _2302_ _2268_ _2303_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_30_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7412_ _3679_ _0414_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_117_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4624_ _1291_ _0737_ _1294_ _1295_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_124_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8392_ _0488_ net1 mod.Data_Mem.F_M.MRAM\[786\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_135_229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_7343_ _3644_ _0380_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4555_ _0653_ mod.Arithmetic.CN.I_in\[58\] mod.Arithmetic.CN.I_in\[59\] _1136_ _1227_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_117_977 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_132_914 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7274_ _3599_ _0356_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4486_ _1153_ _1155_ _1156_ _1157_ _1158_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_116_498 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6225_ _2217_ mod.Data_Mem.F_M.MRAM\[14\]\[3\] mod.Data_Mem.F_M.MRAM\[15\]\[3\] _2319_
+ _2839_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_103_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_1023 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6156_ _2765_ _2770_ _2771_ _2772_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XTAP_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_872 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_894 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5107_ _1563_ _1763_ _1768_ _1773_ _1774_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_97_393 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6087_ _2700_ _2701_ _2703_ _2704_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_45_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5435__A2 _0010_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5038_ _1644_ _1706_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_2706 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2717 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2728 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2739 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6989_ _3405_ mod.Data_Mem.F_M.MRAM\[16\]\[7\] _3428_ _3432_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_55_1130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6902__I _3375_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4946__A1 _1603_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4410__A3 _1082_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_166_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_40_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_1087 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_1128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_154_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8530__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7499__I0 _3645_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_123_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xoutput8 net8 io_out[21] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
Xoutput10 net10 io_out[23] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XFILLER_122_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5253__I _1779_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4477__A3 _0816_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_1156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_682 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_213 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_536 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5831__C1 _2453_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_249 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_964 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_1006 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_32_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8060__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_978 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_82_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_171 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__6139__B1 _2157_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_193 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_121_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_157_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5872__B _2494_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4165__A2 _0840_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5364__S _2025_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4340_ _1009_ _1013_ _1014_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_113_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_119_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5114__A1 _1778_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6259__I _1663_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4271_ _0943_ _0937_ _0944_ _0945_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_67_1089 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5163__I _1816_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6010_ _2413_ _2628_ _2629_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__5665__A2 mod.Data_Mem.F_M.MRAM\[28\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4468__A3 _1140_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_820 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_393 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_503 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7961_ _0187_ net1 mod.Data_Mem.F_M.MRAM\[779\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_82_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6912_ _3249_ mod.Data_Mem.F_M.MRAM\[13\]\[4\] _3381_ _3382_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_36_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_290 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7892_ _0118_ net1 mod.Data_Mem.F_M.MRAM\[25\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__8403__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6843_ _3316_ _3337_ _3344_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_50_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4928__A1 _1594_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5766__C _2376_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6774_ _3295_ _3296_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_50_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3986_ _0640_ mod.Arithmetic.CN.I_in\[64\] _0663_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_8513_ _0017_ net1 mod.Data_Mem.F_M.out_data\[57\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_148_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_22_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5725_ _2068_ _2347_ _2350_ _2168_ _2351_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_50_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8553__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5028__S1 _1651_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8444_ _0540_ net1 mod.Data_Mem.F_M.MRAM\[793\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5656_ _2151_ mod.Data_Mem.F_M.MRAM\[797\]\[2\] _2287_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_136_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4607_ _1162_ _1277_ _1278_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_8375_ _0471_ net1 mod.Data_Mem.F_M.MRAM\[783\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_163_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7553__I _3759_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5587_ _2114_ _2220_ _2224_ _2178_ _0043_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
X_7326_ _3620_ mod.Data_Mem.F_M.MRAM\[770\]\[7\] _3625_ _3633_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_85_1123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_785 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4538_ mod.Arithmetic.CN.I_in\[43\] _1096_ _1210_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_104_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5105__A1 _1769_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7257_ mod.Data_Mem.F_M.MRAM\[31\]\[4\] _3312_ _3590_ _3591_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_85_1178 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4469_ _1087_ _1141_ _1142_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_131_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_104_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6208_ _2779_ _2819_ _2822_ _2692_ _2823_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_7188_ _3549_ _3550_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_58_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_23 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_680 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6139_ mod.Data_Mem.F_M.MRAM\[13\]\[1\] _2751_ _2157_ mod.Data_Mem.F_M.MRAM\[12\]\[1\]
+ _2754_ _2755_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_100_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5801__I _1636_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3204 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3215 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3226 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_3237 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3248 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2503 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3259 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2514 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__4417__I mod.Arithmetic.CN.I_in\[36\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8083__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2525 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2536 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2547 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4092__A1 _0754_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1802 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1813 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2558 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2569 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1824 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1835 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1846 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1857 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_92_1149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1868 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1879 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_31 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_1050 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_167_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_139_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4152__I _0618_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7920__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_155_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4147__A2 _0822_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7463__I _3297_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_123_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6079__I _2295_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_122_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6844__A1 _1955_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5647__A2 _2278_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_122_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_1010 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6807__I _3321_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8426__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_94 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6743__S _3274_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8576__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_753 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5958__I0 mod.Data_Mem.F_M.MRAM\[18\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_639 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4386__A2 mod.Arithmetic.CN.I_in\[20\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7574__S _3773_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5510_ _1779_ _2152_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_6490_ mod.Data_Mem.F_M.MRAM\[12\]\[4\] mod.Data_Mem.F_M.MRAM\[14\]\[4\] mod.Data_Mem.F_M.MRAM\[13\]\[4\]
+ _1870_ _2290_ _2171_ _3095_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_34_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4138__A2 _0709_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_5441_ _2080_ _2077_ _0027_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_145_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5094__S _1746_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7373__I mod.Data_Mem.F_M.MRAM\[773\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4689__A3 _0997_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8160_ mod.Data_Mem.F_M.out_data\[70\] net2 net1 mod.Arithmetic.CN.I_in\[70\] vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_99_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_711 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5372_ mod.Data_Mem.F_M.MRAM\[19\]\[7\] mod.Data_Mem.F_M.MRAM\[18\]\[7\] _1892_ _2034_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_126_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7111_ _3503_ _0289_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_114_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4323_ _0653_ mod.Arithmetic.CN.I_in\[51\] _0997_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__6918__S _3381_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8091_ mod.Data_Mem.F_M.out_data\[1\] net2 net1 mod.Arithmetic.ACTI.x\[1\] vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_99_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5638__A2 _2112_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7042_ _3467_ _0256_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_114_788 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_86_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4254_ _0928_ _0929_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_102_939 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4946__B _1614_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4185_ _0629_ _0853_ _0860_ mod.P3.Res\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_28_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_503 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6438__I1 mod.Data_Mem.F_M.MRAM\[1\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_1059 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_167_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_167_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6063__A2 _2662_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7944_ _0170_ net1 mod.Data_Mem.F_M.MRAM\[789\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_82_344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1109 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_7875_ _0101_ net1 mod.Data_Mem.F_M.MRAM\[24\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_82_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6826_ _3271_ _3332_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_51_753 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7943__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_1160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_797 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6757_ _3285_ _0153_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_23_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_285 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_3969_ _0645_ mod.Arithmetic.CN.I_in\[24\] _0646_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_104_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5708_ _2313_ mod.Data_Mem.F_M.MRAM\[29\]\[6\] _2335_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_12_23 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6688_ _3240_ mod.Data_Mem.F_M.MRAM\[28\]\[1\] _3237_ _3241_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_137_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7315__A2 _3626_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_23 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_8427_ _0523_ net1 mod.Data_Mem.F_M.MRAM\[791\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_100_1109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_5639_ _2265_ _2269_ _2271_ _2272_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_87_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8358_ _0454_ net1 mod.Data_Mem.F_M.MRAM\[781\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__6120__C _2733_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7309_ _3622_ _3623_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_132_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_8289_ _0385_ net1 mod.Data_Mem.F_M.MRAM\[772\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__8449__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5629__A2 _2261_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_714 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_77_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_78_639 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_150_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_609 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_801 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3001 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7626__I0 _3806_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3012 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3023 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_536 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3034 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3045 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2300 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2311 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3056 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_878 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3067 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2322 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3078 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2333 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3089 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2344 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2355 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1610 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2366 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_539 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1621 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1033 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2377 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2388 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1643 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2399 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1654 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1665 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1676 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7554__A2 _3762_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_1200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1687 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1698 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5565__A1 _2070_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5565__B2 _2203_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5907__S _2528_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_154_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6380__I3 mod.Data_Mem.F_M.MRAM\[788\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_1184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5340__I1 mod.Data_Mem.F_M.MRAM\[770\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_801 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5990_ _2079_ _2609_ _2610_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_91_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7966__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_539 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4941_ mod.Data_Mem.F_M.MRAM\[787\]\[0\] mod.Data_Mem.F_M.MRAM\[786\]\[0\] _1609_
+ _1610_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__4851__I0 mod.Data_Mem.F_M.MRAM\[17\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_127_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7660_ mod.Data_Mem.F_M.MRAM\[790\]\[6\] _3824_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4872_ mod.Data_Mem.F_M.src\[0\] _1503_ _1541_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_75_1177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6611_ mod.Data_Mem.F_M.MRAM\[24\]\[1\] _3196_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_20_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7591_ _3785_ _0487_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_60_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6542_ _3083_ mod.Data_Mem.F_M.MRAM\[768\]\[6\] _3145_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_119_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5308__A1 _1942_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6505__B1 _3104_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6473_ _3014_ _3074_ _3078_ _3079_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_134_806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_8212_ _0313_ net1 mod.Data_Mem.F_M.MRAM\[22\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__5859__A2 _2477_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5424_ _1701_ _2081_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_47_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8143_ mod.Data_Mem.F_M.out_data\[53\] net2 net1 mod.Arithmetic.CN.I_in\[53\] vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_114_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5355_ _2012_ _2015_ _2017_ _1822_ _2018_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_82_1126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_160_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4306_ _0891_ mod.Arithmetic.CN.I_in\[35\] _0980_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_8074_ mod.P3.Res\[2\] net2 net1 net5 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_5286_ mod.Data_Mem.F_M.MRAM\[773\]\[5\] mod.Data_Mem.F_M.MRAM\[772\]\[5\] _1612_
+ _1950_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_82_1159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_99_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7025_ _3455_ _0251_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4237_ _0665_ _0846_ _0912_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__4295__A1 _0966_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4168_ _0843_ _0844_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_55_322 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6036__A2 _2156_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_878 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4099_ _0775_ _0776_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_56_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5095__I0 mod.Data_Mem.F_M.MRAM\[773\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6587__A3 _3179_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7927_ _0153_ net1 mod.Data_Mem.F_M.MRAM\[8\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__5795__A1 _2418_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_169_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7858_ _3931_ _0607_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_23_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_572 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6809_ _3323_ _0167_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_169_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8121__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7789_ _3892_ _0578_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_109_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__8271__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_1048 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_2_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_152_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_904 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_574 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_78_469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7989__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_93_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6027__A2 _2641_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_150_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_46_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2130 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2141 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2152 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6306__B _2763_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2163 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2174 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2185 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1440 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1451 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2196 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1462 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1473 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1484 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1495 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_159_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4210__A1 _0881_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5436__I _2069_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_155_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5710__A1 _2071_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5372__S _1892_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_97_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5140_ mod.Data_Mem.F_M.MRAM\[21\]\[3\] mod.Data_Mem.F_M.MRAM\[20\]\[3\] _1510_ _1806_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__5149__S0 _1812_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_393 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5071_ _1737_ _1738_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_81_1181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4022_ _0696_ mod.Arithmetic.I_out\[78\] _0678_ _0698_ _0699_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XFILLER_49_171 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_77_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6018__A2 _2636_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_92_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_539 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8144__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5973_ _2510_ _2591_ _2592_ _2565_ _2593_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__6216__B _2830_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7712_ mod.Data_Mem.F_M.MRAM\[794\]\[0\] _3850_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__8134__D mod.Data_Mem.F_M.out_data\[44\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4924_ _1512_ _1593_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_80_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7643_ _3815_ _0509_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_127_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4855_ _1504_ _1523_ _1524_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__8294__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_159_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7574_ _3747_ mod.Data_Mem.F_M.MRAM\[785\]\[1\] _3773_ _3775_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4786_ mod.Arithmetic.CN.I_in\[15\] _1455_ _1456_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__4201__A1 _0803_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6525_ _2558_ _2598_ _3124_ _3125_ _3128_ _3129_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_146_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_118_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6456_ _3003_ _3055_ _3062_ _3063_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_106_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5407_ _2067_ _2068_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4504__A2 _1062_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_6387_ _2904_ mod.Data_Mem.F_M.MRAM\[783\]\[7\] mod.Data_Mem.F_M.MRAM\[782\]\[7\]
+ _2905_ _2997_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_86_1081 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8126_ mod.Data_Mem.F_M.out_data\[36\] net2 net1 mod.Arithmetic.CN.I_in\[36\] vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_161_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5338_ mod.Data_Mem.F_M.MRAM\[783\]\[6\] _1699_ _2001_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_134_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8057_ _0266_ net1 mod.Data_Mem.F_M.MRAM\[20\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_102_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5269_ _1692_ _1933_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_87_255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7008_ _3443_ _0246_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_75_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6009__A2 _2627_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5068__I0 mod.Data_Mem.F_M.MRAM\[1\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_995 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6804__I1 _3319_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5768__A1 _2382_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5030__B _1697_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6841__S _3340_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7997__RN net2 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4440__A1 mod.Arithmetic.CN.I_in\[52\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_145_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_1014 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6193__A1 _2180_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_138_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5940__A1 _2326_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4743__A2 _1412_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_166_31 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_165_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_125_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_137_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8174__RN net2 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6496__A2 _2559_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_153_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8017__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_1132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_152_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_65_1165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6248__A2 _2224_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_864 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5920__S _2540_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4259__A1 _0907_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_94_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8167__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7048__I1 mod.Data_Mem.F_M.MRAM\[1\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5859__C _2481_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6420__A2 _3025_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7988__RN net2 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4431__A1 _0824_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_572 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1270 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1281 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4982__A2 _1649_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1292 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7646__I mod.Data_Mem.F_M.MRAM\[788\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_1158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4640_ _0695_ _0679_ _1061_ _1311_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__6184__A1 _2070_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6184__B2 _2203_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5231__I0 _1889_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_163_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5931__A1 _2548_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4571_ mod.Arithmetic.CN.I_in\[67\] _1128_ _1243_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__7582__S _3779_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6310_ _1980_ _1981_ _1738_ _2922_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_7290_ _3610_ _3609_ _3611_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_128_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8165__RN net2 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6241_ _1931_ _1857_ _2733_ _2855_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__6487__A2 _3092_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5695__B1 _2323_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_130_116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6172_ _1734_ _1684_ _2775_ _2788_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_124_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_97_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5123_ _1513_ _1790_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6926__S _3391_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_112_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_57_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_85_748 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5054_ _1674_ _1720_ _1721_ _1722_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_38_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5998__A1 _2464_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5998__B2 _2539_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_951 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4005_ mod.Arithmetic.CN.I_in\[18\] _0682_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_38_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4670__A1 _1339_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_995 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5956_ _2531_ _2566_ _2576_ _2577_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__4422__A1 _1091_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4907_ mod.Data_Mem.F_M.MRAM\[774\]\[0\] _1575_ _1576_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5887_ _2506_ mod.Data_Mem.F_M.MRAM\[783\]\[3\] _2507_ _2508_ _2509_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XFILLER_51_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7211__I1 mod.Data_Mem.F_M.MRAM\[2\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4838_ _1506_ _1507_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_7626_ _3806_ mod.Data_Mem.F_M.MRAM\[787\]\[5\] _3801_ _3807_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__6175__A1 _1670_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_575 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5922__A1 _2151_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7557_ _1792_ _3762_ _3764_ _0474_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_4769_ _0624_ _1134_ mod.Arithmetic.CN.I_in\[61\] _1366_ _1439_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_153_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_147_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6508_ _3111_ _3112_ _3113_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_119_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_23 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7488_ _3721_ _0448_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_107_647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_49_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6478__A2 mod.Data_Mem.F_M.MRAM\[769\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6439_ _1619_ _3047_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__8156__RN net2 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5804__I _1903_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_1_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8109_ mod.Data_Mem.F_M.out_data\[19\] net2 net1 mod.Arithmetic.CN.I_in\[19\] vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_0_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5740__S _2358_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5989__A1 _1620_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5989__B2 _2104_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_1084 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_984 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_1103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4661__A1 _1090_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_1125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_43_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6402__A2 mod.Data_Mem.F_M.MRAM\[781\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4413__A1 _1002_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_320 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_169_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_169_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_101_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6166__A1 _1730_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5213__I0 mod.Data_Mem.F_M.MRAM\[1\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_1191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6961__I0 _3399_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4192__A3 _0820_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_1216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8147__RN net2 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6469__A2 mod.Data_Mem.F_M.MRAM\[13\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6713__I0 _3259_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5141__A2 _1601_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6746__S _3279_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_748 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5295__I3 _1958_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_461 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5810_ _2100_ _2434_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_35_678 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_615 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6790_ _3308_ _3309_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_90_784 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5601__B1 _2237_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5741_ _2064_ _2366_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_76_1091 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_128_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_1023 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8460_ _0556_ net1 mod.Data_Mem.F_M.MRAM\[795\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__6157__A1 _2425_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5672_ _2301_ _2213_ _2302_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__6157__B2 _2188_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6213__C _2686_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7411_ mod.Data_Mem.F_M.MRAM\[775\]\[6\] _3679_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4623_ mod.Arithmetic.CN.I_in\[13\] _1189_ _0971_ _1294_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XANTENNA__5904__A1 _2211_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8391_ _0487_ net1 mod.Data_Mem.F_M.MRAM\[785\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__6952__I0 _3386_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7342_ _3615_ mod.Data_Mem.F_M.MRAM\[771\]\[4\] _3643_ _3644_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_128_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4554_ _1225_ _0995_ _1226_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__4949__B _1599_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8332__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8138__RN net2 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7273_ mod.Data_Mem.F_M.MRAM\[5\]\[4\] _3599_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4485_ _1087_ _1141_ _1157_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_89_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6224_ _1931_ _1817_ _2836_ _2837_ _2838_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_106_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6155_ _1910_ _1656_ _2771_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_840 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_1046 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8482__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5106_ _1603_ _1772_ _1651_ _1773_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_895 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6086_ _2702_ _2703_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_57_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5037_ _1702_ _1703_ _1704_ _1705_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_100_878 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2707 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2718 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2729 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_751 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7487__S _3720_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_14_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_1151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5199__A2 _1621_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6988_ _3431_ _0238_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_41_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5939_ _2396_ _2560_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4946__A2 _1613_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6148__A1 _1640_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_1017 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6123__C _2739_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7609_ _3784_ mod.Data_Mem.F_M.MRAM\[786\]\[7\] _3786_ _3796_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_8589_ _0605_ net1 mod.Data_Mem.F_M.MRAM\[9\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_5_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4174__A3 _0849_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8129__RN net2 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7499__I1 mod.Data_Mem.F_M.MRAM\[781\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput9 net9 io_out[22] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XFILLER_123_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6320__A1 _1566_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_1113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_501 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_1168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7120__I0 _3508_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6084__B1 _2165_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_48_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5831__B1 _2451_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5202__C _1699_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_678 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__8205__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6387__A1 _2904_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_71_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_1220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7196__I _3308_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_150 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_161 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_160_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6139__A1 mod.Data_Mem.F_M.MRAM\[13\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__6139__B2 mod.Data_Mem.F_M.MRAM\[12\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_183 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_8_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XPHY_194 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__8355__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_158_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5872__C _1498_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_141_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_114_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4270_ _0865_ _0936_ _0944_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__5380__S _1906_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_79_383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_11_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_67_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7960_ _0186_ net1 mod.Data_Mem.F_M.MRAM\[779\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_54_217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6208__C _2692_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6911_ _3375_ _3381_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_82_548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7891_ _0117_ net1 mod.Data_Mem.F_M.MRAM\[25\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__4009__B mod.Arithmetic.I_out\[72\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6842_ _3343_ _0180_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6378__A1 _2733_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6773_ mod.Data_Mem.F_M.dest\[1\] mod.Data_Mem.F_M.dest\[0\] _3295_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_3985_ _0650_ _0661_ mod.Arithmetic.CN.I_in\[64\] _0662_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XANTENNA__5050__A1 _1714_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5724_ _2280_ _2156_ _2348_ _2349_ _2350_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
X_8512_ _0016_ net1 mod.Data_Mem.F_M.out_data\[56\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_164_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8443_ _0539_ net1 mod.Data_Mem.F_M.MRAM\[793\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5655_ _2091_ _1803_ _2279_ _2286_ _0049_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_50_1050 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_1061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4606_ _1159_ _1196_ _1277_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_129_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8374_ _0470_ net1 mod.Data_Mem.F_M.MRAM\[783\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_50_1072 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6550__A1 _2728_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5586_ mod.Data_Mem.F_M.MRAM\[797\]\[3\] _2179_ _2195_ mod.Data_Mem.F_M.MRAM\[796\]\[3\]
+ _2223_ _2224_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
X_7325_ _3632_ _0374_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_102_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_105_915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4537_ _0654_ mod.Arithmetic.CN.I_in\[44\] _0896_ _0983_ _1209_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XFILLER_2_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7256_ _3584_ _3590_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__5105__A2 mod.Data_Mem.F_M.MRAM\[769\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4468_ _1103_ _1108_ _1140_ _1141_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XANTENNA__7872__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6207_ _2708_ _2820_ _2821_ _2822_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_113_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7187_ _3294_ _3464_ _3335_ _3549_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
X_4399_ _1068_ _1069_ _1071_ _1072_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_113_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6138_ _2752_ _2753_ _2754_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_320 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6066__B1 mod.Data_Mem.F_M.MRAM\[783\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3205 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3216 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6069_ _2685_ _2686_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_3227 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8228__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3238 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3249 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2504 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2515 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2526 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2537 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2548 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1803 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2559 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1814 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6369__A1 _2869_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1825 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1836 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_497 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1847 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1858 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8378__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1869 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_158_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5529__I _1915_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7169__I0 _3539_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_1062 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6916__I0 _3256_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_154_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6541__A1 _2091_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5344__A2 _2006_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4147__A3 _0669_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_123_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_1208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6844__A2 _3337_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_110_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4855__A1 _1504_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_153_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_49_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_504 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4607__A1 _1162_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5280__A1 _1941_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_44_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_765 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5958__I1 mod.Data_Mem.F_M.MRAM\[19\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4343__I mod.Arithmetic.CN.I_in\[59\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_73_1050 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_160_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_41_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_1045 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_73_1094 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6907__I0 _3243_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_1089 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5440_ _2072_ _2074_ _2076_ _0026_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XANTENNA__6532__A1 _2061_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7895__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5371_ mod.Data_Mem.F_M.MRAM\[21\]\[7\] mod.Data_Mem.F_M.MRAM\[20\]\[7\] _1890_ _2033_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_126_561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7590__S _3779_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7110_ _3450_ mod.Data_Mem.F_M.MRAM\[3\]\[1\] _3501_ _3503_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_113_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4322_ _0891_ mod.Arithmetic.CN.I_in\[50\] _0838_ _0996_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
X_8090_ mod.Data_Mem.F_M.out_data\[0\] net2 net1 mod.Arithmetic.ACTI.x\[0\] vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_99_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_113_233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5099__A1 _1708_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6296__B1 mod.Data_Mem.F_M.MRAM\[782\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7041_ _3445_ mod.Data_Mem.F_M.MRAM\[1\]\[0\] _3466_ _3467_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4253_ mod.Arithmetic.CN.I_in\[50\] _0928_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_113_288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4184_ _0748_ _0855_ _0857_ _0859_ _0628_ _0860_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_132_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7943_ _0169_ net1 mod.Data_Mem.F_M.MRAM\[789\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__5271__A1 _1933_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8520__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7874_ _0100_ net1 mod.Data_Mem.F_M.MRAM\[24\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_63_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_169_929 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_50_220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6825_ _3331_ _0175_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_51_765 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7765__S _3878_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4253__I mod.Arithmetic.CN.I_in\[50\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6756_ mod.Data_Mem.F_M.MRAM\[8\]\[1\] _3285_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_50_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_1172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3968_ _0641_ _0645_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_5707_ _2334_ _0053_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_6687_ _3239_ _3240_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_136_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8426_ _0522_ net1 mod.Data_Mem.F_M.MRAM\[791\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__6523__A1 _2315_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5638_ _2270_ _2112_ _2271_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_163_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_152_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_8357_ _0453_ net1 mod.Data_Mem.F_M.MRAM\[781\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__5084__I _1524_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5569_ _2184_ _2207_ _2208_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_117_572 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7308_ _3332_ _3604_ _3446_ _3622_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_132_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_8288_ _0384_ net1 mod.Data_Mem.F_M.MRAM\[772\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_105_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7239_ _3580_ _0340_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_104_277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8050__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7005__S _3440_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4837__A1 _1499_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4301__A3 _0974_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_651 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_504 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3002 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3013 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3024 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3035 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3046 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2301 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3057 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2312 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3068 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2323 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2334 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3079 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1600 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_163_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2345 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2356 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_710 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1611 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2367 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1622 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2378 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1633 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2389 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1644 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_148_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_1655 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1666 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_169_31 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_159_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1677 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_169_42 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_787 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1688 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_169_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_1212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_155_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6514__A1 _2475_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6311__C _2078_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_1196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_607 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4828__A1 _1493_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_748 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8543__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_846 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_643 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4940_ _1509_ _1609_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_45_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4851__I1 mod.Data_Mem.F_M.MRAM\[16\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_91_197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_32_220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4871_ mod.Data_Mem.F_M.MRAM\[5\]\[0\] mod.Data_Mem.F_M.MRAM\[4\]\[0\] _1514_ _1540_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_2890 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4073__I _0710_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6610_ _3195_ _0096_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_7590_ _3784_ mod.Data_Mem.F_M.MRAM\[785\]\[7\] _3779_ _3785_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_32_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6541_ _2091_ _2622_ _3143_ _3144_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_9_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6472_ _3021_ _2527_ _2524_ _3009_ _3077_ _3078_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XANTENNA__6505__A1 _2611_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5308__A2 mod.Data_Mem.F_M.MRAM\[0\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6505__B2 _2211_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_145_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_118_358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8211_ _0312_ net1 mod.Data_Mem.F_M.MRAM\[22\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5423_ _2080_ _2077_ _0011_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_134_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6929__S _3391_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__8073__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5354_ _1704_ _2016_ _2017_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_8142_ mod.Data_Mem.F_M.out_data\[52\] net2 net1 mod.Arithmetic.CN.I_in\[52\] vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_114_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4305_ _0895_ _0899_ _0979_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_141_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8073_ mod.P3.Res\[1\] net2 net1 net4 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_5285_ _1927_ _1930_ _1948_ _1949_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_99_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5867__I0 mod.Data_Mem.F_M.MRAM\[14\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7024_ _3454_ mod.Data_Mem.F_M.MRAM\[18\]\[3\] _3448_ _3455_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4236_ _0664_ _0846_ _0911_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__5492__A1 _2135_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4295__A2 _0968_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4248__I _0922_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_971 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4167_ mod.Arithmetic.CN.F_in\[0\] _0843_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_95_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7910__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4098_ mod.Arithmetic.ACTI.x\[3\] _0775_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_82_153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5095__I1 mod.Data_Mem.F_M.MRAM\[772\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7926_ _0152_ net1 mod.Data_Mem.F_M.MRAM\[8\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_55_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_1201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7857_ mod.Data_Mem.F_M.MRAM\[9\]\[7\] _3931_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5079__I _1518_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_169_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_142_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6808_ mod.Data_Mem.F_M.MRAM\[799\]\[7\] _3322_ _3313_ _3323_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_23_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_168_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7788_ _3306_ mod.Data_Mem.F_M.MRAM\[798\]\[2\] _3889_ _3892_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_11_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4755__B1 _1213_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_1021 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6739_ _3240_ mod.Data_Mem.F_M.MRAM\[0\]\[1\] _3274_ _3276_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_20_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_137_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8416__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7544__I0 _3729_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_1016 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4507__B1 _1064_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8409_ _0505_ net1 mod.Data_Mem.F_M.MRAM\[788\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__6839__S _3340_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5743__S _1515_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5970__C _2572_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_155_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8566__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_78_426 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_31 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4286__A2 _0808_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_610 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3997__I mod.Arithmetic.CN.I_in\[23\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5235__B2 _1897_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_1009 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2120 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2131 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_34_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2142 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2153 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2164 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2175 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1430 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2186 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1441 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2197 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1452 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1463 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1474 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1485 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1496 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5717__I _1691_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8096__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_116_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5710__A2 _2148_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5149__S1 _1814_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4496__C _1072_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_746 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7933__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5070_ _1606_ _1737_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_85_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4021_ mod.Arithmetic.I_out\[77\] _0698_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_81_1193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_429 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_930 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5972_ mod.Data_Mem.F_M.MRAM\[14\]\[5\] mod.Data_Mem.F_M.MRAM\[15\]\[5\] _2528_ _2592_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__5777__A2 _1548_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_646 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6216__C _2374_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7711_ _3849_ _0543_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4923_ _1583_ _1591_ _1558_ _1592_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__8439__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7642_ mod.Data_Mem.F_M.MRAM\[788\]\[5\] _3815_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4854_ _1522_ _1492_ _1523_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__7774__I0 _3778_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4785_ _1288_ _0735_ _1455_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_7573_ _3774_ _0480_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4201__A2 _0875_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4531__I _1202_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6524_ _2500_ _2602_ _3127_ _3128_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__8589__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6455_ _3056_ _3057_ _3061_ _3014_ _3062_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_162_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5406_ _2066_ _2067_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6386_ mod.Data_Mem.F_M.MRAM\[13\]\[7\] _1538_ _2201_ mod.Data_Mem.F_M.MRAM\[12\]\[7\]
+ _2995_ _2996_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_115_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5337_ _1986_ _1992_ _1993_ _1999_ _1899_ _2000_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
X_8125_ mod.Data_Mem.F_M.out_data\[35\] net2 net1 mod.Arithmetic.CN.I_in\[35\] vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_88_713 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_130_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8056_ _0265_ net1 mod.Data_Mem.F_M.MRAM\[20\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5268_ _1890_ _1932_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_76_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7007_ _3403_ mod.Data_Mem.F_M.MRAM\[17\]\[6\] _3440_ _3443_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4219_ _0820_ _0826_ _0894_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_69_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5199_ mod.Data_Mem.F_M.MRAM\[799\]\[3\] _1621_ _1625_ _1865_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_21_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5068__I1 mod.Data_Mem.F_M.MRAM\[0\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_985 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5768__A2 _2384_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_1140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7909_ _0135_ net1 mod.Data_Mem.F_M.MRAM\[28\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_71_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_1004 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__4440__A2 _0997_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_1075 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7765__I0 _3293_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6193__A2 _1735_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_109_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_164_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_125_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7956__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_152_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_3_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_746 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_843 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_1177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4259__A2 _0927_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5456__A1 _2081_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_90_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4616__I mod.Arithmetic.CN.I_in\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_163_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6008__I0 mod.Data_Mem.F_M.MRAM\[770\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6831__I _3336_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1260 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1271 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_124_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1282 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1293 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6184__A2 mod.Data_Mem.F_M.MRAM\[14\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6052__B _2666_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5447__I _1522_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5231__I1 _1891_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4195__A1 _0638_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_156_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4570_ mod.Arithmetic.CN.I_in\[66\] _1129_ _0634_ _0775_ _1242_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XFILLER_7_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_155_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6240_ _2160_ _1853_ _2854_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5144__B1 _1808_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5695__A1 _2082_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6278__I _2228_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5695__B2 _2306_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6171_ _1645_ _1680_ _2787_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_69_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5122_ _1714_ mod.Data_Mem.F_M.MRAM\[787\]\[2\] _1788_ _1789_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_97_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8111__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_278 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5053_ _1507_ _1721_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_69_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5998__A2 _2615_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__4954__C _1622_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4004_ mod.Arithmetic.I_out\[75\] _0681_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_84_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_974 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_65_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8261__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_432 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_52_145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5955_ _2410_ _2570_ _2573_ _2575_ _2576_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_40_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4906_ _1574_ _1575_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_5886_ _2209_ _2508_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_61_690 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7625_ _3315_ _3806_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4837_ _1499_ _1505_ _1506_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_21_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6175__A2 _2778_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7979__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7556_ _3612_ _3762_ _3764_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_5_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5922__A2 _1919_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4768_ mod.Arithmetic.ACTI.x\[7\] _1436_ _1437_ _1438_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_88_1111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_146_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6507_ _3049_ _2323_ _2500_ _2543_ _2541_ _2568_ _3112_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XANTENNA__4981__I0 mod.Data_Mem.F_M.MRAM\[1\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4699_ _0891_ mod.Arithmetic.CN.I_in\[69\] _1370_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_7487_ _3718_ mod.Data_Mem.F_M.MRAM\[781\]\[0\] _3720_ _3721_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__5135__B1 _1760_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_1188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6438_ mod.Data_Mem.F_M.MRAM\[0\]\[1\] mod.Data_Mem.F_M.MRAM\[1\]\[1\] _2512_ _3046_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_161_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6369_ _2869_ _2978_ _2979_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_8108_ mod.Data_Mem.F_M.out_data\[18\] net2 net1 mod.Arithmetic.CN.I_in\[18\] vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_103_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_716 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5438__A1 _2089_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8039_ _0248_ net1 mod.Data_Mem.F_M.MRAM\[18\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_75_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4110__A1 _0781_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4110__B2 _0786_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_646 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_432 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__5610__A1 _2228_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4413__A2 _1022_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8092__RN net2 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_24_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5267__I _1695_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6166__A2 _1711_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5213__I1 mod.Data_Mem.F_M.MRAM\[0\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_536 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6961__I1 _1870_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_165_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_6_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_137_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_819 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6713__I1 mod.Data_Mem.F_M.MRAM\[28\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8134__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5677__A1 _2135_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_532 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5730__I _2354_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8284__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_568 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4652__A2 _1322_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_432 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_50_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5601__A1 _2225_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5378__S _1814_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4404__A2 _1075_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5601__B2 _2178_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5740_ mod.Data_Mem.F_M.MRAM\[18\]\[0\] mod.Data_Mem.F_M.MRAM\[19\]\[0\] _2358_ _2365_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_76_1081 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_690 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1090 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_89_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5671_ _1692_ _2301_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_50_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7410_ _3678_ _0413_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4622_ _1291_ _1292_ _1293_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_8390_ _0486_ net1 mod.Data_Mem.F_M.MRAM\[785\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__6952__I1 mod.Data_Mem.F_M.MRAM\[15\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_773 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7341_ _3635_ _3643_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_4553_ mod.Arithmetic.CN.I_in\[52\] _1225_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_116_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7272_ _3598_ _0355_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4484_ _1087_ _1141_ _1156_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__5668__A1 _2068_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6223_ _2714_ _2685_ _2837_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_143_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_44_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6154_ _1751_ _1659_ _2770_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_830 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_83_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_852 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_513 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4891__A2 _1552_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6736__I _3273_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5105_ _1769_ mod.Data_Mem.F_M.MRAM\[769\]\[2\] _1771_ _1772_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6085_ _2209_ _2201_ _2702_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_100_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_248 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5140__I0 mod.Data_Mem.F_M.MRAM\[21\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5036_ _1573_ _1704_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_2708 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_122_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_39_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_66_771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5840__A1 _2085_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2719 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_66_782 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_730 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6987_ _3403_ mod.Data_Mem.F_M.MRAM\[16\]\[6\] _3428_ _3431_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_53_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8074__RN net2 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5288__S _1951_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_80_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8007__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5938_ mod.Data_Mem.F_M.MRAM\[16\]\[4\] mod.Data_Mem.F_M.MRAM\[17\]\[4\] _2189_ _2559_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_34_690 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5869_ _2124_ _2454_ _2367_ _2490_ _2491_ _2170_ _2492_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XANTENNA__4159__A1 _0830_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7608_ _3795_ _0494_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4920__S _1588_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8588_ _0604_ net1 mod.Data_Mem.F_M.MRAM\[9\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_126_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8157__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_166_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_147_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_7539_ _3725_ _1901_ _3752_ _3753_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_107_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5815__I _2422_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6847__S _3336_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_116_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__6320__A2 _1936_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_163_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_513 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_102_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7120__I1 mod.Data_Mem.F_M.MRAM\[3\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_546 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6084__A1 _2081_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6084__B2 _1620_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7820__A2 _3908_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5831__A1 _2449_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_730 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_752 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_914 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6387__A2 mod.Data_Mem.F_M.MRAM\[783\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4398__A1 _0871_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_34_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_162 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6139__A2 _2751_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__5926__S _2339_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_184 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__5898__A1 _2118_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_154_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_1203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4322__A1 _0891_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_39_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5822__A1 _2416_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6910_ _3380_ _0211_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_7890_ _0116_ net1 mod.Data_Mem.F_M.MRAM\[25\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_63_752 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6841_ _3249_ mod.Data_Mem.F_M.MRAM\[769\]\[4\] _3340_ _3343_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_165_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_51_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6291__I _2059_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_1198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5586__B1 _2195_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6772_ _3229_ _3294_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_51_969 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3984_ mod.Arithmetic.ACTI.x\[0\] _0661_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__6224__C _2837_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8511_ net187 net1 mod.Data_Mem.F_M.out_data\[71\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5723_ _1932_ mod.Data_Mem.F_M.MRAM\[796\]\[7\] _2217_ _2349_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__5836__S _2152_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8442_ _0538_ net1 mod.Data_Mem.F_M.MRAM\[793\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_31_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5654_ _2068_ _2285_ _2286_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_148_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4605_ _1154_ _1274_ _1275_ _1276_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_8373_ _0469_ net1 mod.Data_Mem.F_M.MRAM\[783\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__5635__I _2267_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6550__A2 mod.Data_Mem.F_M.MRAM\[1\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5585_ _2221_ _2222_ _2223_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_129_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_1084 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7324_ _3618_ mod.Data_Mem.F_M.MRAM\[770\]\[6\] _3625_ _3632_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4536_ _0651_ mod.Arithmetic.CN.I_in\[45\] _1208_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_85_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7255_ _3589_ _0347_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_131_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4467_ _1121_ _1122_ _1139_ _1140_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_89_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4313__A1 _0982_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6206_ _1730_ _1767_ _2821_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_7186_ _3548_ _0319_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4398_ _0871_ _1064_ _1070_ _1071_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_86_800 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_14 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6137_ _2009_ mod.Data_Mem.F_M.MRAM\[14\]\[1\] mod.Data_Mem.F_M.MRAM\[15\]\[1\] _1968_
+ _2753_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XTAP_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_682 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_855 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6066__A1 _2517_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6066__B2 _2567_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3206 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_85_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3217 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6068_ _1676_ _2375_ _1495_ _2685_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_86_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3228 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_1191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5813__A1 _2321_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3239 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2505 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5019_ mod.Data_Mem.F_M.MRAM\[788\]\[1\] _1687_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_2516 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2527 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2538 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1804 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2549 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1815 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_785 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1826 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_936 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1837 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1848 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1859 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_13_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7318__A1 _3555_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7169__I1 mod.Data_Mem.F_M.MRAM\[12\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__6526__C1 _2606_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6916__I1 mod.Data_Mem.F_M.MRAM\[13\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_710 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5545__I _1533_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6541__A2 _2622_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_765 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_123_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_162_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_107_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5481__S _1845_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4304__A1 _0901_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4304__B2 _0907_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_150_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_682 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4097__S _0746_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_535 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_546 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6057__A1 _2288_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_85 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7201__S _3553_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8322__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_33_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_72_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_788 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_1084 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4791__A1 mod.Arithmetic.CN.I_in\[23\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6517__C1 _2580_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8472__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_158_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_118_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6907__I1 mod.Data_Mem.F_M.MRAM\[13\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6532__A2 mod.Data_Mem.F_M.MRAM\[1\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4543__A1 mod.Arithmetic.CN.I_in\[35\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5370_ mod.Data_Mem.F_M.MRAM\[23\]\[7\] mod.Data_Mem.F_M.MRAM\[22\]\[7\] _1588_ _2032_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_160_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_154_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4321_ _0654_ _0928_ mod.Arithmetic.CN.I_in\[51\] _0995_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_113_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6296__A1 _2144_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7040_ _3465_ _3466_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__6296__B2 _2267_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5343__I0 _2002_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4252_ _0910_ _0921_ _0926_ _0927_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_99_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_1180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_1033 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4183_ _0748_ _0858_ _0795_ _0859_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_68_844 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6048__A1 _2560_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7942_ _0168_ net1 mod.Data_Mem.F_M.MRAM\[789\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_94_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5271__A2 _1934_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7873_ _0099_ net1 mod.Data_Mem.F_M.MRAM\[24\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__6235__B _2718_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6824_ mod.Data_Mem.F_M.MRAM\[789\]\[7\] _3331_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_50_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6220__A1 _2832_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6755_ _3284_ _0152_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_52_1113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3967_ _0643_ mod.Arithmetic.CN.I_in\[16\] _0644_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_91_1184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5706_ _2082_ _2329_ _2333_ _2306_ _2334_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_164_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6686_ net4 _3239_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_8425_ _0521_ net1 mod.Data_Mem.F_M.MRAM\[791\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5637_ _1811_ _2270_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__6523__A2 _1955_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8201__RN net2 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4534__A1 _1203_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8356_ _0452_ net1 mod.Data_Mem.F_M.MRAM\[781\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_128_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5568_ _2159_ _2206_ _1631_ _2207_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_89_1080 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_29 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7307_ _3621_ _0367_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4519_ _0724_ _0707_ _0971_ _1191_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_8287_ _0383_ net1 mod.Data_Mem.F_M.MRAM\[771\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_144_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5499_ _1879_ mod.Data_Mem.F_M.MRAM\[30\]\[5\] _2143_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_104_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6287__B2 _2899_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7238_ _3533_ mod.Data_Mem.F_M.MRAM\[30\]\[4\] _3579_ _3580_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__5334__I0 mod.Data_Mem.F_M.MRAM\[17\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4837__A2 _1505_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7169_ _3539_ mod.Data_Mem.F_M.MRAM\[12\]\[7\] _3534_ _3540_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_58_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_150_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6039__A1 _2288_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3003 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8345__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3014 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3025 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6834__I0 _3240_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_160_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3036 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2302 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_3047 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7021__S _3448_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3058 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2313 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3069 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2324 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2335 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2346 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1601 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2357 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1612 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_571 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1623 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2368 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_722 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_891 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2379 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1634 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_42_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1645 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8495__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1656 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6211__A1 _1706_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1678 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1689 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6514__A2 _1971_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_142_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_64_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_111_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_49_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6450__A1 _2696_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_91_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2880 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4870_ _1538_ _1539_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_2891 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6202__A1 _2681_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7250__I0 _1632_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7862__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6540_ _2619_ mod.Data_Mem.F_M.MRAM\[780\]\[6\] _3142_ _2170_ _3143_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_146_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_159_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_71_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6471_ _2422_ _3075_ _3076_ _3077_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XANTENNA__6505__A2 _2547_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8210_ _0311_ net1 mod.Data_Mem.F_M.MRAM\[12\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__8218__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4516__A1 _0824_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5422_ _2079_ _2080_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_86_1220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_161_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_893 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_8141_ mod.Data_Mem.F_M.out_data\[51\] net2 net1 mod.Arithmetic.CN.I_in\[51\] vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_5353_ mod.Data_Mem.F_M.MRAM\[785\]\[6\] mod.Data_Mem.F_M.MRAM\[784\]\[6\] _1580_
+ _2016_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_126_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5913__I _1726_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5316__I0 mod.Data_Mem.F_M.MRAM\[19\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4304_ _0901_ _0902_ _0934_ _0977_ _0907_ _0978_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai32_1
XFILLER_88_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8072_ mod.P3.Res\[0\] net2 net1 net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_114_576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5284_ _1551_ _1939_ _1947_ _1948_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__8368__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7023_ _3245_ _3454_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5867__I1 mod.Data_Mem.F_M.MRAM\[15\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5134__B _1800_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4235_ _0841_ _0908_ _0909_ _0910_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_101_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5492__A2 mod.Data_Mem.F_M.MRAM\[30\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4166_ _0807_ mod.Arithmetic.CN.I_in\[65\] _0842_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_55_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_782 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4097_ mod.Arithmetic.CN.I_in\[11\] _0721_ _0746_ _0774_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_55_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7925_ _0151_ net1 mod.Data_Mem.F_M.MRAM\[0\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_82_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6992__A2 _3371_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7776__S _3883_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_7856_ _3930_ _0606_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_24_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_169_749 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6807_ _3321_ _3322_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_7787_ _3891_ _0577_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4999_ _1657_ _1660_ _1662_ _1666_ _1616_ _1667_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XANTENNA__4755__A1 mod.Arithmetic.CN.I_in\[37\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6738_ _3275_ _0144_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_104_1000 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_165_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6669_ mod.Data_Mem.F_M.MRAM\[27\]\[6\] _3225_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_104_1055 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7544__I1 mod.Data_Mem.F_M.MRAM\[783\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8408_ _0504_ net1 mod.Data_Mem.F_M.MRAM\[788\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__4507__A1 _0632_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_152_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_104_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_830 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_8339_ _0435_ net1 mod.Data_Mem.F_M.MRAM\[778\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_151_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_120_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_150_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_63_1094 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_1113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_74_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_1157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_62_806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6432__A1 _1965_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2110 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7480__I0 _3618_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2121 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7885__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2132 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2143 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2154 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2165 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1420 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2176 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1431 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1442 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_64_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2187 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2198 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_14_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1453 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_159_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1464 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1475 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1497 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4746__A1 mod.Arithmetic.CN.I_in\[69\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6322__C _1866_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_155_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_115_307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8510__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_108_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5733__I _1681_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4020_ mod.Arithmetic.CN.I_in\[23\] _0677_ _0697_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_96_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_38_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5971_ mod.Data_Mem.F_M.MRAM\[2\]\[5\] mod.Data_Mem.F_M.MRAM\[3\]\[5\] _2540_ _2591_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_18_571 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7710_ mod.Data_Mem.F_M.MRAM\[793\]\[7\] _3849_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_80_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4922_ _1585_ _1589_ _1590_ _1591_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_61_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7223__I0 _3537_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7641_ _3814_ _0508_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4037__I0 _0687_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4853_ _1521_ _1522_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__7774__I1 mod.Data_Mem.F_M.MRAM\[797\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8040__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7572_ _3771_ mod.Data_Mem.F_M.MRAM\[785\]\[0\] _3773_ _3774_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4784_ _0743_ _1294_ _1453_ _1454_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_147_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6523_ _2315_ _1955_ _2406_ _3126_ _3127_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_101_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6454_ _2503_ _2478_ _3059_ _2568_ _3060_ _2477_ _3061_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_133_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8190__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5405_ _1724_ _2065_ _2066_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__5162__A1 _1826_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6385_ _1565_ _2994_ _2995_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_133_148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_1072 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8124_ mod.Data_Mem.F_M.out_data\[34\] net2 net1 mod.Arithmetic.CN.I_in\[34\] vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_5336_ _1888_ _1998_ _1633_ _1999_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_138_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8055_ _0264_ net1 mod.Data_Mem.F_M.MRAM\[20\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_47_1078 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_87_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_130_855 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5267_ _1695_ _1931_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_69_961 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7006_ _3442_ _0245_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_60_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4218_ mod.Arithmetic.CN.I_in\[34\] _0893_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_87_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5198_ mod.Data_Mem.F_M.MRAM\[783\]\[3\] _1863_ _1864_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_29_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4149_ _0824_ mod.Arithmetic.CN.I_in\[48\] _0668_ _0825_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_56_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_997 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4208__B _0882_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_1010 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7908_ _0134_ net1 mod.Data_Mem.F_M.MRAM\[28\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_58_1152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7839_ _3169_ _3921_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_70_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_54_1049 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7765__I1 mod.Data_Mem.F_M.MRAM\[797\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8533__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_153_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_119_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4878__B _1533_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_117_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_714 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_121_822 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4259__A3 _0933_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5456__A2 _2104_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_717 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_87_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5502__B _2084_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_942 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_93_249 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_677 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8063__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_91 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7205__I0 _3539_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6008__I1 mod.Data_Mem.F_M.MRAM\[771\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1250 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1261 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1272 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_91_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_1283 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1294 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4719__A1 _1273_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5231__I2 _1893_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5392__A1 _2012_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7900__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_116_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5144__B2 _1809_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_1212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5695__A2 _2318_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6170_ _2196_ _1689_ _2739_ _2786_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_112_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_69_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5121_ _1715_ _1787_ _1788_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_123_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_85_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5052_ _1700_ _1705_ _1712_ _1719_ _1720_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_111_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_739 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4003_ mod.Arithmetic.CN.I_in\[19\] _0680_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__8406__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_603 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5131__C _1558_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_168_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5954_ _2506_ _1870_ _2075_ _2574_ _2575_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_4905_ _1573_ _1574_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_52_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_1216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8556__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_680 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5885_ _2266_ mod.Data_Mem.F_M.MRAM\[782\]\[3\] _2507_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__6243__B _2743_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7624_ _1919_ _3804_ _3805_ _0500_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_33_393 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4836_ _1501_ _1504_ _1505_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_21_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_166_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7555_ _1678_ _3762_ _3763_ _0473_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_4767_ mod.Arithmetic.CN.I_in\[68\] _1377_ _1422_ mod.Arithmetic.ACTI.x\[5\] _1437_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XFILLER_53_1093 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6506_ _2107_ _3111_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_135_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_107_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7486_ _3719_ _3720_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_88_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4698_ _0620_ _1367_ _1368_ _1369_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_134_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_107_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_1156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5135__A1 _1729_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_162_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6437_ _2312_ _2459_ _3044_ _3026_ _3045_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__5135__B2 _1670_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6368_ _2974_ _2975_ _2976_ _2977_ _2978_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_103_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_103_822 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8107_ mod.Data_Mem.F_M.out_data\[17\] net2 net1 mod.Arithmetic.CN.I_in\[17\] vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_0_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5319_ _1551_ _1982_ _1508_ _1983_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_102_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6299_ _2232_ _2237_ _2908_ _2911_ _1964_ _2759_ _2912_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_8038_ _0247_ net1 mod.Data_Mem.F_M.MRAM\[17\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_103_888 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_60_1020 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_739 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_611 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4110__A2 _0780_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8086__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_56_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_147_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_1149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_147_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5997__I0 mod.Data_Mem.F_M.MRAM\[784\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_322 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA_output10_I net10 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_71_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5548__I _2187_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_169_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_169_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__7923__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_588 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_1171 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5126__A1 _1715_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_152_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_133_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8429__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_971 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_982 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5232__B _1633_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_430 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_75_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8579__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_62_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5601__A2 _2232_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4404__A3 _1076_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_15_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5458__I _2106_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1080 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1091 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5670_ _2270_ _2127_ _2300_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_148_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4621_ _0731_ _1191_ _1292_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_11_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7340_ _3642_ _0379_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_117_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_11_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4552_ _1118_ _1119_ _1223_ _1224_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_128_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_144_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6289__I _1543_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7271_ mod.Data_Mem.F_M.MRAM\[5\]\[3\] _3598_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4483_ _1047_ _1084_ _1155_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_104_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5668__A2 _2298_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6222_ _1734_ _1819_ _2836_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_83_1020 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4876__B1 _1531_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6153_ _2759_ _2764_ _2768_ _2769_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XTAP_820 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_48_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_1015 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7114__S _3501_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_853 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_717 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_503 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5104_ _1708_ _1770_ _1771_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_98_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_864 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_875 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6084_ _2081_ _1497_ _2165_ _1620_ _1965_ _2701_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_112_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_897 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7290__A1 _3610_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6093__A2 _2708_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5035_ mod.Data_Mem.F_M.MRAM\[775\]\[1\] mod.Data_Mem.F_M.MRAM\[774\]\[1\] _1692_
+ _1703_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__5140__I1 mod.Data_Mem.F_M.MRAM\[20\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_964 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_100_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_38_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2709 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6986_ _3430_ _0237_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_54_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_606 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7946__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_797 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5937_ _2402_ _2558_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_53_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7784__S _3889_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5868_ mod.Data_Mem.F_M.MRAM\[16\]\[2\] mod.Data_Mem.F_M.MRAM\[17\]\[2\] _2152_ _2491_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_55_1177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_167_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7607_ _3782_ mod.Data_Mem.F_M.MRAM\[786\]\[6\] _3786_ _3795_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4819_ _1267_ _1485_ _1486_ _1487_ _1488_ mod.P3.Res\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__oai32_1
XANTENNA__4159__A2 _0834_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8587_ _0603_ net1 mod.Data_Mem.F_M.MRAM\[9\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5799_ _2422_ _2423_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_7538_ _3744_ _3752_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_107_402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7469_ _3709_ _0441_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_134_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_107_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_820 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_27_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_153_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7024__S _3448_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_48_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_674 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6084__A2 _1497_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5831__A2 _2450_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5595__A1 mod.Data_Mem.F_M.MRAM\[29\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4398__A2 _1064_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5595__B2 mod.Data_Mem.F_M.MRAM\[28\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5278__I _1514_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_130 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_152 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_163 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_169_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_185 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__8101__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_157_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4910__I _1578_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8194__191 net191 vdd vss gf180mcu_fd_sc_mcu7t5v0__tieh
XANTENNA__5898__A2 _2505_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_1004 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8251__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_119_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4322__A2 mod.Arithmetic.CN.I_in\[50\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_1215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_503 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7969__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6840_ _3342_ _0179_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_62_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_904 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6771_ _3292_ _3293_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_3983_ _0659_ _0660_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_90_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8510_ net188 net1 mod.Data_Mem.F_M.out_data\[70\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_50_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5722_ _2281_ mod.Data_Mem.F_M.MRAM\[797\]\[7\] _2348_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_149_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8441_ _0537_ net1 mod.Data_Mem.F_M.MRAM\[793\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__5338__A1 mod.Data_Mem.F_M.MRAM\[783\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5653_ _2280_ _2121_ _2282_ _2284_ _2285_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XANTENNA__6521__B _2596_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4820__I mod.Data_Mem.F_M.src\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4604_ _1158_ _1258_ _1275_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_8372_ _0468_ net1 mod.Data_Mem.F_M.MRAM\[783\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5584_ _2138_ mod.Data_Mem.F_M.MRAM\[799\]\[3\] mod.Data_Mem.F_M.MRAM\[798\]\[3\]
+ _2088_ _2222_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_7_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7323_ _3631_ _0373_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_117_755 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_1096 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4535_ _1206_ _1207_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_85_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7254_ mod.Data_Mem.F_M.MRAM\[31\]\[3\] _3555_ _3585_ _3589_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4466_ _1133_ _1138_ _1139_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_116_287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_427 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6205_ _1706_ _1772_ _2820_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_120_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7185_ mod.Data_Mem.F_M.MRAM\[22\]\[7\] _3548_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5651__I _1779_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4397_ _0843_ mod.Arithmetic.CN.I_in\[28\] _1070_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_112_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6136_ _1564_ _2752_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_536 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_569 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6067_ _2682_ _2683_ _2684_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_3207 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3218 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3229 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5018_ _1594_ _1686_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_2506 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2517 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2528 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2539 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1805 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1816 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_572 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1827 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1838 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5577__A1 _2214_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1849 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8124__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6969_ _3419_ _0231_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_42_23 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7318__A2 _3623_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_981 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_158_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6526__B1 _3060_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6526__C2 _3107_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8274__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_166_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_108_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_755 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5501__A1 _2144_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5561__I _1538_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_801 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_131_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6057__A2 mod.Data_Mem.F_M.MRAM\[4\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4905__I _1573_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7557__A2 _3762_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5568__A1 _2159_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_981 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6517__B1 _3050_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6517__C2 _2496_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_160_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4543__A2 _1091_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4320_ _0922_ _0660_ _0840_ _0994_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_114_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_99_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4251_ _0923_ _0924_ _0925_ _0926_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XANTENNA__5343__I1 _2003_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_113_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_1192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4182_ _0763_ _0764_ _0858_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_122_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_110_931 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA_input1_I io_in[8] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_1007 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_1089 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7941_ _0167_ net1 mod.Data_Mem.F_M.MRAM\[799\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__8147__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_167_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_48_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7872_ _0098_ net1 mod.Data_Mem.F_M.MRAM\[24\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_36_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6008__S _2275_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_169_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6823_ _3330_ _0174_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5559__A1 _2196_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8297__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6220__A2 _2833_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6754_ mod.Data_Mem.F_M.MRAM\[8\]\[0\] _3284_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_17_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3966_ _0642_ _0643_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_91_1152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5705_ _2316_ _2142_ _2330_ _2332_ _2333_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XANTENNA__4782__A2 _1451_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6685_ _3238_ _0128_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_52_1169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8424_ _0520_ net1 mod.Data_Mem.F_M.MRAM\[791\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5636_ _2266_ mod.Data_Mem.F_M.MRAM\[28\]\[0\] _2268_ _2269_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_148_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_128_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_164_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8355_ _0451_ net1 mod.Data_Mem.F_M.MRAM\[781\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__5731__A1 _2187_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5567_ mod.Data_Mem.F_M.MRAM\[29\]\[2\] _2200_ _2202_ mod.Data_Mem.F_M.MRAM\[28\]\[2\]
+ _2205_ _2206_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_2
XFILLER_89_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7306_ _3620_ mod.Data_Mem.F_M.MRAM\[768\]\[7\] _3608_ _3621_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4518_ _1189_ _1190_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_8286_ _0382_ net1 mod.Data_Mem.F_M.MRAM\[771\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_2_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5498_ _1778_ mod.Data_Mem.F_M.MRAM\[798\]\[5\] _2141_ _2142_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_7237_ _3573_ _3579_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__6287__A2 _2885_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6477__I _2189_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5334__I1 mod.Data_Mem.F_M.MRAM\[16\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4449_ _1007_ _1015_ _1016_ _1105_ _1122_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XFILLER_120_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_160_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7168_ _3258_ _3539_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_98_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_942 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6119_ mod.Data_Mem.F_M.MRAM\[23\]\[0\] mod.Data_Mem.F_M.MRAM\[22\]\[0\] _1782_ _2736_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_19_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_59_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7099_ _3496_ _0284_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_74_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3004 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_101_986 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3015 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3026 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_539 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3037 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3048 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2303 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3059 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2314 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2325 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2336 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2347 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1602 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2358 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1613 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2369 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1624 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1085 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1646 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1058 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_169_11 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1657 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1668 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6211__A2 _1794_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1679 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_149_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_168_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5970__A1 _2587_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5556__I _1639_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_167_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5722__A1 _2281_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4525__A2 _1162_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_154_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_108_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_155_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_123_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_322 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_290 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_675 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_91 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_1103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2870 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2881 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2892 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_1169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7250__I1 _3303_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4213__A1 _0825_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5961__A1 _2475_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6071__B _1729_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_119_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6470_ _2275_ mod.Data_Mem.F_M.MRAM\[12\]\[3\] _3076_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_5421_ _2078_ _2079_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_146_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8195__RN net2 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5713__A1 _2339_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4516__A2 _0731_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_127_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_160_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_500 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8140_ mod.Data_Mem.F_M.out_data\[50\] net2 net1 mod.Arithmetic.CN.I_in\[50\] vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_5352_ _1933_ _2013_ _2014_ _2015_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_99_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4303_ _0927_ _0933_ _0977_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_8071_ mod.DMen_reg net2 net1 mod.DMen_reg2 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_99_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5283_ _1805_ _1944_ _1946_ _1947_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__5316__I1 mod.Data_Mem.F_M.MRAM\[18\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_717 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7022_ _3453_ _0250_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_87_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4234_ _0619_ _0661_ mod.Arithmetic.CN.I_in\[64\] _0847_ _0909_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_114_17 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4165_ _0659_ _0840_ _0841_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__7122__S _3506_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_461 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4096_ _0754_ _0766_ _0767_ _0773_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_82_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6961__S _3414_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7924_ _0150_ net1 mod.Data_Mem.F_M.MRAM\[0\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_70_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4452__A1 _0614_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7855_ mod.Data_Mem.F_M.MRAM\[9\]\[6\] _3930_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6806_ net10 _3321_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_23_255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4998_ _1664_ _1665_ _1666_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_51_575 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7786_ _3303_ mod.Data_Mem.F_M.MRAM\[798\]\[1\] _3889_ _3891_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_11_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6737_ _3228_ mod.Data_Mem.F_M.MRAM\[0\]\[0\] _3274_ _3275_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_108_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3949_ _0626_ mod.DM_en vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5952__A1 _2062_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4755__A2 _1423_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_1023 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6668_ _3224_ _0125_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_128_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_149_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8407_ _0503_ net1 mod.Data_Mem.F_M.MRAM\[787\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5619_ _2233_ mod.Data_Mem.F_M.MRAM\[799\]\[7\] mod.Data_Mem.F_M.MRAM\[798\]\[7\]
+ _2229_ _2253_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_165_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6752__I0 _3259_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5704__A1 _2331_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_1029 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6599_ mod.Data_Mem.F_M.MRAM\[11\]\[3\] _3190_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_136_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8338_ _0434_ net1 mod.Data_Mem.F_M.MRAM\[778\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_105_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_105_533 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8312__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8269_ _0365_ net1 mod.Data_Mem.F_M.MRAM\[768\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_78_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6000__I _1778_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_675 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8462__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_1125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_101_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_100_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_859 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6432__A2 _3039_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_1169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2100 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7480__I1 mod.Data_Mem.F_M.MRAM\[780\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8110__RN net2 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2111 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2122 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4443__A1 _0915_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2133 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2144 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1410 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2155 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2166 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1421 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2177 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1432 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2188 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1443 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2199 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1465 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6196__A1 _1751_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1476 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1487 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1498 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_35_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_1180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5943__A1 _2558_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4746__A2 _1376_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8177__RN net2 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6743__I0 _3246_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_465 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_155_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_89_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_97_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_69_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6120__A1 _1505_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6120__B2 _1575_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_96_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_1162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4682__A1 mod.Arithmetic.CN.I_in\[61\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_77_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8101__RN net2 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5970_ _2587_ mod.Data_Mem.F_M.MRAM\[5\]\[5\] _2589_ _2572_ _2590_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_92_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4921_ _1561_ _1590_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_45_380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_391 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7223__I1 mod.Data_Mem.F_M.MRAM\[2\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7640_ mod.Data_Mem.F_M.MRAM\[788\]\[4\] _3814_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4852_ mod.Data_Mem.F_M.src\[0\] _1521_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__6187__A1 _2687_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4037__I1 _0683_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_7571_ _3772_ _3773_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_21_759 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5934__A1 _2379_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4783_ _0743_ _1190_ _1188_ _1453_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_165_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_159_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_140_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6522_ _2321_ mod.Data_Mem.F_M.MRAM\[768\]\[5\] _3126_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__8335__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8168__RN net2 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6453_ _2499_ _3060_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_147_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7117__S _3506_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5404_ _2064_ _1553_ _2065_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_161_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_680 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6384_ _2134_ mod.Data_Mem.F_M.MRAM\[15\]\[7\] mod.Data_Mem.F_M.MRAM\[14\]\[7\] _2216_
+ _2994_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__5162__A2 _1827_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8123_ mod.Data_Mem.F_M.out_data\[33\] net2 net1 mod.Arithmetic.CN.I_in\[33\] vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_5335_ _1994_ _1995_ _1996_ _1997_ _1844_ _1882_ _1998_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_87_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8485__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_1016 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_8054_ _0263_ net1 mod.Data_Mem.F_M.MRAM\[1\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5266_ mod.Data_Mem.F_M.MRAM\[799\]\[5\] _1599_ _1930_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_87_225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_536 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7005_ _3416_ mod.Data_Mem.F_M.MRAM\[17\]\[5\] _3440_ _3442_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4217_ _0891_ mod.Arithmetic.CN.I_in\[34\] _0892_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_130_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_68_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5197_ _1557_ _1863_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4673__A1 _1334_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_56_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4148_ _0620_ _0824_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__7611__A1 _3296_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4079_ _0754_ _0708_ _0721_ _0722_ _0756_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__4425__A1 _0619_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5622__B1 _2255_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7907_ _0133_ net1 mod.Data_Mem.F_M.MRAM\[28\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_55_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7586__I _3318_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_1164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6178__A1 _2319_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7838_ _3920_ _0610_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_51_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6178__B2 _2311_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_169_569 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_157_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7769_ _3306_ mod.Data_Mem.F_M.MRAM\[797\]\[2\] _3878_ _3881_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_50_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_166_23 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8159__RN net2 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_606 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_3_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5055__B _1722_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_1157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6102__A1 _2186_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4113__B1 _0789_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_47_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4664__A1 _1202_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8524__182 net182 vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_86_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8208__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4416__A1 _0982_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_497 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_90_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_391 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8532__D _0036_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_163_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7205__I1 mod.Data_Mem.F_M.MRAM\[29\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1240 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1251 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6169__A1 _2186_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_575 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1262 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1284 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8358__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1295 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5916__A1 _2428_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6964__I0 _3416_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_147_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5231__I3 _1895_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5392__A2 _2051_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_680 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5144__A2 _1645_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5120_ mod.Data_Mem.F_M.MRAM\[786\]\[2\] _1787_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_97_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7141__I0 _3460_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7841__A1 _0610_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5051_ _1713_ _1718_ _1651_ _1719_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_112_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_46_1090 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_66_910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4002_ _0678_ _0679_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_84_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_751 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4095__I _0768_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_26_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_66_987 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4407__A1 _0715_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_1017 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5953_ _2266_ mod.Data_Mem.F_M.MRAM\[14\]\[4\] _2574_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_81_968 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6524__B _3127_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5919__I _1783_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4823__I mod.Data_Mem.F_M.src\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4904_ _1572_ _1573_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_21_501 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5884_ _2319_ _2506_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_139_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7623_ _3312_ _3804_ _3805_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_4835_ _1502_ _1503_ _1504_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__5855__S _2398_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7554_ _3610_ _3762_ _3763_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_4766_ _1422_ mod.Arithmetic.ACTI.x\[7\] _1436_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_140_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_119_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6505_ _2611_ _2547_ _3104_ _2211_ _3109_ _3110_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_88_1113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_1004 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7485_ _3634_ _3371_ _3387_ _3719_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_4697_ _1134_ _1250_ _1366_ _1368_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or3_1
XFILLER_107_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6436_ _2071_ _3042_ _3043_ _3044_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_88_1168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5135__A2 _1627_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__7875__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6367_ _1834_ _2028_ _2873_ _2977_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_115_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5318_ _1978_ _1979_ _1980_ _1981_ _1527_ _1795_ _1982_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_8106_ mod.Data_Mem.F_M.out_data\[16\] net2 net1 mod.Arithmetic.CN.I_in\[16\] vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_88_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7132__I0 _3452_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6298_ mod.Data_Mem.F_M.MRAM\[781\]\[4\] _2751_ _2157_ mod.Data_Mem.F_M.MRAM\[780\]\[4\]
+ _2910_ _2911_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_102_344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8037_ _0246_ net1 mod.Data_Mem.F_M.MRAM\[17\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5249_ _1503_ _1914_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_88_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_1054 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6399__A1 _3004_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_1117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7310__S _3623_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_497 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8500__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_312 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__7199__I0 _3533_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_323 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_52_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_24_383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_12_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_169_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5765__S _1951_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_71_1183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5564__I _2096_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_153_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_126_948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_69_1090 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6395__I _2698_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8030__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4637__A1 _0633_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_74_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_710 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8180__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4643__I mod.Arithmetic.CN.I_in\[30\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_1081 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_163_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_1015 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_37_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_31_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1092 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6011__B1 _2625_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4620_ _0828_ _1289_ _1290_ _1291_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__6562__A1 _2385_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7898__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4551_ _0929_ _1113_ _1115_ _1116_ _1112_ _1223_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
X_7270_ _3597_ _0354_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4482_ _0988_ _1083_ _1153_ _1154_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_132_907 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6221_ mod.Data_Mem.F_M.MRAM\[1\]\[3\] mod.Data_Mem.F_M.MRAM\[2\]\[3\] mod.Data_Mem.F_M.MRAM\[3\]\[3\]
+ mod.Data_Mem.F_M.MRAM\[4\]\[3\] _2588_ _2449_ _2835_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_98_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4876__A1 mod.Data_Mem.F_M.MRAM\[3\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_1190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_1092 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6152_ _2765_ _2766_ _2767_ _2768_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XTAP_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7114__I0 _3454_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_832 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_843 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5103_ mod.Data_Mem.F_M.MRAM\[768\]\[2\] _1770_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_97_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6083_ _1802_ _2697_ _2699_ _2700_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_100_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_876 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4628__A1 _1185_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_887 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_898 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5034_ mod.Data_Mem.F_M.MRAM\[773\]\[1\] mod.Data_Mem.F_M.MRAM\[772\]\[1\] _1701_
+ _1702_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_111_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8523__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_924 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7130__S _3513_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6985_ _3416_ mod.Data_Mem.F_M.MRAM\[16\]\[5\] _3428_ _3430_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_53_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_54_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4553__I mod.Arithmetic.CN.I_in\[52\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5936_ _2366_ _2556_ _2100_ _2449_ _2557_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_80_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_1161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_34_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_5867_ mod.Data_Mem.F_M.MRAM\[14\]\[2\] mod.Data_Mem.F_M.MRAM\[15\]\[2\] _2452_ _2490_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_51_1009 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_166_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7606_ _3794_ _0493_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_21_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4818_ _0673_ _0674_ mod.Arithmetic.I_out\[79\] _0675_ _1488_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_1
XANTENNA__6553__A1 _2343_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8586_ _0602_ net1 mod.Data_Mem.F_M.MRAM\[9\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_21_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5798_ _1596_ _2422_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_5_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7537_ _3751_ _0467_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4749_ _0623_ mod.Arithmetic.CN.I_in\[70\] _1379_ _1419_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_135_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_119_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6305__A1 _1655_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_162_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5739__S0 _1714_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7468_ _3638_ mod.Data_Mem.F_M.MRAM\[780\]\[1\] _3707_ _3709_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_134_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6419_ _2626_ _3027_ _3028_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_7399_ mod.Data_Mem.F_M.MRAM\[775\]\[0\] _3673_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__8053__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_88_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6148__C _2763_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5292__A1 _1875_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6943__I _3255_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_968 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5044__A1 _1706_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_1212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_120 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_71_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_131 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_158_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_142 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_153 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_169_185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_9_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_197 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_8_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_1016 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_607 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_158_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_981 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7215__S _3562_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4322__A3 _0838_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__8546__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7014__I _3447_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6058__C _2572_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_751 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5283__A1 _1805_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_1123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_0 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_90_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5586__A2 _2179_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3982_ _0635_ mod.Arithmetic.CN.I_in\[56\] _0659_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6770_ net3 _3292_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_5721_ _2312_ _2154_ _2344_ _2346_ _2347_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_94_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_148_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8440_ _0536_ net1 mod.Data_Mem.F_M.MRAM\[793\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__5338__A2 _1699_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6535__A1 _3060_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5652_ _2283_ mod.Data_Mem.F_M.MRAM\[28\]\[1\] _2217_ _2284_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__6535__B2 _3020_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_164_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_50_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_1042 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4603_ _1158_ _1258_ _1274_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_5583_ _1549_ _2221_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_8371_ _0467_ net1 mod.Data_Mem.F_M.MRAM\[783\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_117_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8076__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7322_ _3569_ mod.Data_Mem.F_M.MRAM\[770\]\[5\] _3625_ _3631_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4534_ _1203_ _1098_ _1206_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_144_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7253_ _3588_ _0346_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_85_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4465_ _0923_ _1135_ _1137_ _1138_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_137_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6204_ _1566_ _1761_ _1762_ _1555_ _2819_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_131_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7184_ _3547_ _0318_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_131_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4396_ _0615_ _0958_ _1063_ _1055_ _1069_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XANTENNA__6249__B _2862_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_651 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_640 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6135_ _1538_ _2751_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_113_984 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6964__S _3414_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_651 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_133_16 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_526 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7913__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6066_ _2517_ mod.Data_Mem.F_M.MRAM\[782\]\[0\] mod.Data_Mem.F_M.MRAM\[783\]\[0\]
+ _2567_ _2683_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_100_645 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4992__B _1614_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3208 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_1171 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5274__A1 _1645_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3219 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5017_ _1518_ _1685_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_38_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_710 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2507 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2518 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_66_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_96_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2529 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5600__C _2236_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_765 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1806 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5026__A1 _1691_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1817 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1828 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1839 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6968_ _3405_ mod.Data_Mem.F_M.MRAM\[15\]\[7\] _3414_ _3419_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_53_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5919_ _1783_ _2540_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_6899_ mod.Data_Mem.F_M.dest\[4\] _3372_ _3373_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_50_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_167_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_1054 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6526__A1 _2508_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5329__A2 _1991_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8419__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7574__I0 _3747_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6526__B2 _2605_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8569_ _0073_ net1 mod.Data_Mem.F_M.out_data\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_107_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7326__I0 _3620_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_163_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8569__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6938__I _3390_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_150_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5501__A2 mod.Data_Mem.F_M.MRAM\[31\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8077__D mod.P3.Res\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_526 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_49_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_87 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6673__I net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5289__I _1579_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5568__A2 _2206_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_1020 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_164_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_41_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8099__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4921__I _1561_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6517__A1 _3049_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7565__I0 _3729_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6517__B2 _2578_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_157_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_146_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_118_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_153_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4250_ _0637_ _0922_ _0924_ _0925_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__7936__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4181_ _0856_ _0857_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4059__A2 _0730_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5256__A1 _1918_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7940_ _0166_ net1 mod.Data_Mem.F_M.MRAM\[799\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_48_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6516__C _2434_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7871_ _0097_ net1 mod.Data_Mem.F_M.MRAM\[24\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_169_1081 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_871 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_169_1092 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6822_ mod.Data_Mem.F_M.MRAM\[789\]\[6\] _3330_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_90_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_90_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6753_ _3283_ _0151_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_50_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3965_ _0641_ _0642_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_149_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4831__I mod.Data_Mem.F_M.src\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_1164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5704_ _2331_ mod.Data_Mem.F_M.MRAM\[796\]\[5\] _2088_ _2332_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__6024__S _2528_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6684_ _3228_ mod.Data_Mem.F_M.MRAM\[28\]\[0\] _3237_ _3238_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_8423_ _0519_ net1 mod.Data_Mem.F_M.MRAM\[790\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__3990__A1 _0662_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5635_ _2267_ _2268_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5863__S _1954_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_8354_ _0450_ net1 mod.Data_Mem.F_M.MRAM\[781\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_145_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5731__A2 _1499_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5566_ _1664_ _2204_ _2205_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_105_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7305_ _3321_ _3620_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4517_ mod.Arithmetic.CN.I_in\[12\] _1189_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_8285_ _0381_ net1 mod.Data_Mem.F_M.MRAM\[771\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5497_ _1686_ mod.Data_Mem.F_M.MRAM\[799\]\[5\] _2141_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_132_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7236_ _3578_ _0339_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_104_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4448_ _1111_ _1120_ _1121_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__5495__A1 _2138_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_59_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7167_ _3538_ _0310_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4379_ _0687_ _0804_ _1050_ _1051_ _1052_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_99_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6118_ _2373_ _2687_ _2730_ _2731_ _2734_ _2735_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XTAP_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_643 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_7098_ mod.Data_Mem.F_M.MRAM\[23\]\[4\] _3496_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_85_131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7589__I _3321_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5247__A1 _1552_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_86_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3005 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3016 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3027 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6049_ _1612_ mod.Data_Mem.F_M.MRAM\[19\]\[7\] _2667_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XTAP_3038 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3049 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2304 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1020 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2315 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_96_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2326 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2337 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2348 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1603 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1614 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2359 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1625 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8241__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1636 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7795__I0 _3806_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1647 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1658 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_169_23 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1669 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_1204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4741__I _1338_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5970__A2 mod.Data_Mem.F_M.MRAM\[5\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_128_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8391__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3981__A1 _0636_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7959__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5722__A2 mod.Data_Mem.F_M.MRAM\[797\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_151_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_68_1188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5486__A1 _1799_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_2_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7227__A2 _3464_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_816 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6038__I0 mod.Data_Mem.F_M.MRAM\[770\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_166_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_584 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_893 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2860 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_32_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2871 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_32_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7786__I0 _3303_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2882 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2893 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4213__A2 _0849_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_430 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6779__S _3300_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5420_ _1489_ _2078_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_127_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5713__A2 mod.Data_Mem.F_M.MRAM\[796\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_1200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5351_ _1903_ mod.Data_Mem.F_M.MRAM\[786\]\[6\] _2014_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_57_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_47_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4302_ _0952_ _0975_ _0976_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_99_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5282_ _1826_ _1945_ _1946_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_8070_ _0279_ net1 mod.Data_Mem.F_M.MRAM\[21\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__8114__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7021_ _3452_ mod.Data_Mem.F_M.MRAM\[18\]\[2\] _3448_ _3453_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4233_ _0662_ _0847_ _0908_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_102_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4164_ _0617_ mod.Arithmetic.CN.I_in\[57\] _0840_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_114_29 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4826__I mod.Data_Mem.F_M.src\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4095_ _0768_ _0772_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_82_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8264__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7923_ _0149_ net1 mod.Data_Mem.F_M.MRAM\[0\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_71_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_819 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4452__A2 mod.Arithmetic.CN.I_in\[68\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7854_ _3929_ _0605_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_64_893 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_690 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_169_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6805_ _3320_ _0166_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_51_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5657__I _1609_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7785_ _3890_ _0576_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4997_ mod.Data_Mem.F_M.MRAM\[21\]\[1\] mod.Data_Mem.F_M.MRAM\[20\]\[1\] _1636_ _1665_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_23_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6736_ _3273_ _3274_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_3948_ mod.P1.instr_reg\[17\] _0625_ _0626_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_6667_ mod.Data_Mem.F_M.MRAM\[27\]\[5\] _3224_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_8406_ _0502_ net1 mod.Data_Mem.F_M.MRAM\[787\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_30_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5618_ mod.Data_Mem.F_M.MRAM\[29\]\[7\] _2086_ _1639_ mod.Data_Mem.F_M.MRAM\[28\]\[7\]
+ _2251_ _2252_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XFILLER_164_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5704__A2 mod.Data_Mem.F_M.MRAM\[796\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6598_ _3189_ _0090_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6752__I1 mod.Data_Mem.F_M.MRAM\[0\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_8337_ _0433_ net1 mod.Data_Mem.F_M.MRAM\[778\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5549_ _1790_ _2189_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_2_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_8268_ _0364_ net1 mod.Data_Mem.F_M.MRAM\[768\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_105_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_160_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7219_ _3568_ _0332_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_8199_ _0084_ net2 net1 mod.I_addr\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_48_23 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4140__A1 _0621_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6437__B _3044_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2101 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2112 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6283__I3 mod.Data_Mem.F_M.MRAM\[788\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2123 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4443__A2 mod.Arithmetic.CN.I_in\[52\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2134 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5640__A1 _2084_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_161_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6951__I _3408_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2145 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1400 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4672__S _1342_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2156 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1411 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2167 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_64_77 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_746 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1433 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2178 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2189 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1444 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1455 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6196__A2 _1747_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1466 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6172__B _2775_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1477 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1488 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_168_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1499 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5943__A2 _2559_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_1192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3954__A1 _0622_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_1056 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_70_1078 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_167_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6743__I1 mod.Data_Mem.F_M.MRAM\[0\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8137__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_157_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_7_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5251__S0 _1829_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4420__B _0826_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4847__S _1515_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_150_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8287__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7223__S _3567_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6347__B _2739_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_985 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_1185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_462 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_93_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_540 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4920_ mod.Data_Mem.F_M.MRAM\[769\]\[0\] mod.Data_Mem.F_M.MRAM\[768\]\[0\] _1588_
+ _1589_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_33_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7759__I0 _3782_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2690 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4851_ mod.Data_Mem.F_M.MRAM\[17\]\[0\] mod.Data_Mem.F_M.MRAM\[16\]\[0\] _1519_ _1520_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__6187__A2 _2801_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_166_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_61_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4198__A1 _0807_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7570_ _3705_ _3335_ _3758_ _3772_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_4782_ _1447_ _1451_ _1452_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_14_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_158_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_140_1213 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6521_ _2567_ mod.Data_Mem.F_M.MRAM\[780\]\[5\] _2596_ _3125_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_6452_ _2345_ _1770_ _3058_ _3059_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_146_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5403_ _1501_ _2064_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6383_ _2979_ _2982_ _2989_ _2992_ _2993_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__4330__B _1003_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8122_ mod.Data_Mem.F_M.out_data\[32\] net2 net1 mod.Arithmetic.CN.I_in\[32\] vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_115_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5334_ mod.Data_Mem.F_M.MRAM\[17\]\[6\] mod.Data_Mem.F_M.MRAM\[16\]\[6\] _1894_ _1997_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_130_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_142_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8053_ _0262_ net1 mod.Data_Mem.F_M.MRAM\[1\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_87_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5265_ _1929_ _0004_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_134_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_930 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__4984__C _1651_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7004_ _3441_ _0244_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4216_ _0653_ _0891_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_102_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5196_ _1552_ _1825_ _1861_ _1862_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_56_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_782 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4147_ _0821_ _0822_ _0669_ _0823_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_68_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_793 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_56_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_95_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4078_ _0750_ _0751_ _0708_ _0754_ _0755_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XANTENNA__5622__A1 _2225_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4425__A2 mod.Arithmetic.CN.I_in\[41\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5622__B2 _2177_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6771__I _3292_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7906_ _0132_ net1 mod.Data_Mem.F_M.MRAM\[28\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_58_1121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_690 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7837_ _3913_ _3915_ _3919_ _3920_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_52_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_145_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6178__A2 mod.Data_Mem.F_M.MRAM\[783\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_169_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_51_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7768_ _3880_ _0569_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6719_ mod.Data_Mem.F_M.MRAM\[10\]\[2\] _3263_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_7_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7699_ _3843_ _0537_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_149_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_165_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5689__A1 _2312_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5336__B _1633_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7107__I _3500_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4361__A1 _0781_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_161_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6946__I _3258_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_1169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6102__A2 _1582_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7043__S _3466_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4113__A1 _0786_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4113__B2 mod.Arithmetic.ACTI.x\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4664__A2 mod.Arithmetic.CN.I_in\[45\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5861__A1 _2416_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_793 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8095__RN net2 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5613__A1 _1940_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4416__A2 _1088_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6681__I _3234_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_163_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1230 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1252 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6413__I0 mod.Data_Mem.F_M.MRAM\[0\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1263 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_513 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1274 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1285 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1296 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_129_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_42_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6964__I1 mod.Data_Mem.F_M.MRAM\[15\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7218__S _3567_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_155_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7017__I _3239_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_1203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_640 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_124_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5760__I _1840_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_151_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7141__I1 mod.Data_Mem.F_M.MRAM\[19\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5050_ _1714_ mod.Data_Mem.F_M.MRAM\[769\]\[1\] _1717_ _1718_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_38_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4001_ mod.Arithmetic.CN.I_in\[21\] _0678_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_78_771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_782 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_1061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_168_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_38_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_53_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5604__A1 mod.Data_Mem.F_M.MRAM\[29\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5604__B2 mod.Data_Mem.F_M.MRAM\[28\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5952_ _2062_ mod.Data_Mem.F_M.MRAM\[5\]\[4\] _2571_ _2572_ _2573_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_18_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4903_ _1571_ _1572_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__8302__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5883_ _2423_ _2131_ _2498_ _2504_ _2505_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_7622_ _3801_ _3804_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_21_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4834_ mod.Data_Mem.F_M.src\[1\] _1503_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_159_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_7553_ _3759_ _3762_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_14_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4765_ _1359_ _1360_ _1434_ _1358_ _1435_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__7128__S _3513_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6504_ _3105_ _3108_ _2474_ _3109_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__6032__S _2331_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8452__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7484_ _3292_ _3718_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_147_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4696_ _1134_ _1250_ _1366_ _1367_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_119_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6435_ _2417_ mod.Data_Mem.F_M.MRAM\[13\]\[1\] _3043_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_161_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6332__A2 _2935_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6366_ _1941_ _2027_ _2976_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_1_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8105_ mod.Data_Mem.F_M.out_data\[15\] net2 net1 mod.Arithmetic.CN.I_in\[15\] vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_143_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5317_ mod.Data_Mem.F_M.MRAM\[17\]\[5\] mod.Data_Mem.F_M.MRAM\[16\]\[5\] _1568_ _1981_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_88_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7132__I1 mod.Data_Mem.F_M.MRAM\[19\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6297_ _2752_ _2909_ _2910_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_103_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8036_ _0245_ net1 mod.Data_Mem.F_M.MRAM\[17\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_76_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_568 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5248_ _1672_ _1913_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_130_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_25_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_1180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_57_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5843__A1 _2417_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_68_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5179_ _1578_ _1845_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_57_977 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6399__A2 _3007_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8077__RN net2 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_785 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_796 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_1129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_690 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__7199__I1 mod.Data_Mem.F_M.MRAM\[29\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_335 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_129_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6020__A1 _2185_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_71_1151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6450__B _2382_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_71_1195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4582__A1 _1249_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_67_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4334__A1 _0640_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_106_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6087__A1 _2700_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7823__A2 _3908_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_48_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4637__A2 _0958_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8325__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5598__B1 mod.Data_Mem.F_M.MRAM\[798\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_788 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1071 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8475__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1082 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1093 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6011__A1 _2379_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6011__B2 _2626_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4022__B1 _0678_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6562__A2 mod.Data_Mem.F_M.MRAM\[768\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_398 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4573__A1 _1125_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4550_ _1121_ _1220_ _1221_ _1222_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_128_264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6787__S _3300_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4481_ _1047_ _1084_ _1153_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_6220_ _2832_ _2833_ _2834_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5373__I0 mod.Data_Mem.F_M.MRAM\[17\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5522__B1 mod.Data_Mem.F_M.MRAM\[31\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_125_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4876__A2 _1539_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5704__B _2088_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6151_ _2180_ _1649_ _2767_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_800 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5490__I _2134_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7114__I1 mod.Data_Mem.F_M.MRAM\[3\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_822 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_643 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_844 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5102_ _1701_ _1769_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_97_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_855 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6082_ mod.Data_Mem.F_M.MRAM\[13\]\[0\] _2087_ _2212_ mod.Data_Mem.F_M.MRAM\[12\]\[0\]
+ _2698_ _2699_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_112_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4628__A2 _1093_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_888 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5033_ _1676_ _1701_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_66_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_988 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_796 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4834__I mod.Data_Mem.F_M.src\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6984_ _3429_ _0236_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_1133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_65_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_755 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6250__A1 _2212_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5935_ mod.Data_Mem.F_M.MRAM\[18\]\[4\] mod.Data_Mem.F_M.MRAM\[19\]\[4\] _2301_ _2556_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_22_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_34_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5866_ _2447_ _2488_ _2489_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_90_1037 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6002__A1 _2620_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7050__I0 _3456_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7605_ _3754_ mod.Data_Mem.F_M.MRAM\[786\]\[5\] _3787_ _3794_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_21_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4817_ _0797_ _0672_ _1487_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_8585_ _0601_ net1 mod.Data_Mem.F_M.MRAM\[9\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__8231__RN net2 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6553__A2 mod.Data_Mem.F_M.MRAM\[13\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5797_ _2110_ _2420_ _2421_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_108_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7536_ _3711_ mod.Data_Mem.F_M.MRAM\[783\]\[3\] _3745_ _3751_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__4564__A1 _1234_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4748_ _1414_ _1415_ _1417_ _1418_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_135_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_119_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7467_ _3708_ _0440_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_107_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6305__A2 _1974_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4679_ _1224_ _1232_ _1350_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__5739__S1 _1756_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4316__A1 _0988_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7992__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5364__I0 mod.Data_Mem.F_M.MRAM\[3\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6418_ _3026_ _2272_ _2365_ _3006_ _2361_ _2672_ _3027_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_116_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7398_ _3672_ _0407_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_134_278 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_162_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6349_ _2869_ _2959_ _2960_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_88_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_131_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__8348__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4619__A2 mod.Arithmetic.CN.I_in\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8019_ _0228_ net1 mod.Data_Mem.F_M.MRAM\[15\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_48_229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_538 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_730 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_432 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5292__A2 mod.Data_Mem.F_M.MRAM\[768\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_722 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_17_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8498__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6241__A1 _1931_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5044__A2 _1711_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_132 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_71_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_169_142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_12_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_52_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_143 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_160_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_154 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__7041__I0 _3445_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_165 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_8_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_187 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_169_197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_40_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4555__A1 _0653_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_166_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_21_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4307__A1 _0893_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4307__B2 mod.Arithmetic.CN.I_in\[33\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_79_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5807__A1 _2428_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7231__S _3574_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6480__A1 _3031_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_1168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_1179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_917 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_165_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_1 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_63_788 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_574 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7865__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3981_ _0636_ mod.Arithmetic.CN.I_in\[48\] _0658_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_44_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5720_ _2345_ mod.Data_Mem.F_M.MRAM\[28\]\[7\] _2280_ _2346_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__4794__A1 _1423_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5651_ _1779_ _2283_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_87_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6535__A2 _2643_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_1021 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4602_ _0625_ _0735_ _1190_ _1079_ _1273_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
X_8370_ _0466_ net1 mod.Data_Mem.F_M.MRAM\[783\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_30_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5582_ _2211_ _2212_ _2219_ _2220_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_7321_ _3630_ _0372_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_50_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4533_ _1203_ _1099_ _1204_ _1095_ _1205_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_156_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_102_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6310__S _1738_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7252_ mod.Data_Mem.F_M.MRAM\[31\]\[2\] _3306_ _3585_ _3588_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_116_256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4464_ _0923_ _1019_ _1136_ _1137_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_144_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6203_ _2810_ _2817_ _2818_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__4829__I _1497_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7183_ mod.Data_Mem.F_M.MRAM\[22\]\[6\] _3547_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4395_ _0956_ _1059_ _1068_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XTAP_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6134_ _2685_ _2750_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_674 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6065_ _2681_ _2682_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3209 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5274__A2 _1937_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6471__A1 _2422_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_1183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5016_ _1675_ mod.Data_Mem.F_M.MRAM\[787\]\[1\] _1683_ _1684_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_85_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_26_402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_1213 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2508 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6980__S _3423_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2519 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_81_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1807 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1818 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1829 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6967_ _3418_ _0230_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_53_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5918_ _2402_ _2539_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_107_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6898_ mod.Data_Mem.F_M.dest\[2\] _3372_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_166_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5849_ _2439_ _2125_ _2469_ _2403_ _2471_ _2472_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XANTENNA__6526__A2 _2333_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8020__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4537__A1 _0654_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8568_ _0072_ net1 mod.Data_Mem.F_M.out_data\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_108_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_154_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_148_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_713 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7519_ _3740_ _0460_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__7326__I1 mod.Data_Mem.F_M.MRAM\[770\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8499_ _0003_ net1 mod.Data_Mem.F_M.out_data\[75\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_107_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8170__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_1072 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_1_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_153_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6837__I0 _3243_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_67_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7888__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4863__I2 _1516_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6214__A1 _1898_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_1010 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4776__A1 _1300_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_158_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_60_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_1054 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_160_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6517__A2 _2329_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_1049 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7565__I1 mod.Data_Mem.F_M.MRAM\[784\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4528__A1 _1108_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5725__B1 _2350_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8513__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_5_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_749 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4180_ _0797_ mod.P2.Rout_reg\[1\] _0856_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_68_836 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5256__A2 _1919_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7870_ _0096_ net1 mod.Data_Mem.F_M.MRAM\[24\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__6205__A1 _1706_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6821_ _3329_ _0173_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_23_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_1110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8043__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6752_ _3259_ mod.Data_Mem.F_M.MRAM\[0\]\[7\] _3279_ _3283_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__4767__A1 mod.Arithmetic.CN.I_in\[68\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3964_ _0640_ _0641_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__7005__I0 _3416_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_148_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5703_ _1581_ _2331_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_6683_ _3236_ _3237_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_91_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6508__A2 _3112_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8422_ _0518_ net1 mod.Data_Mem.F_M.MRAM\[790\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_164_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5634_ _1493_ _2267_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__3990__A2 _0666_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8193__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5192__A1 _1844_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8353_ _0449_ net1 mod.Data_Mem.F_M.MRAM\[781\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5565_ _2070_ mod.Data_Mem.F_M.MRAM\[30\]\[2\] mod.Data_Mem.F_M.MRAM\[31\]\[2\] _2203_
+ _2204_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_163_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7304_ _3619_ _0366_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4516_ _0824_ _0731_ _1188_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_8284_ _0380_ net1 mod.Data_Mem.F_M.MRAM\[771\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_160_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5496_ _2119_ _2137_ _2140_ _2133_ _0036_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
X_7235_ _3531_ mod.Data_Mem.F_M.MRAM\[30\]\[3\] _3574_ _3578_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4447_ _1118_ _1119_ _1120_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_104_237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_63_1201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5495__A2 mod.Data_Mem.F_M.MRAM\[798\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_1212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7166_ _3537_ mod.Data_Mem.F_M.MRAM\[12\]\[6\] _3534_ _3538_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_99_983 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4378_ _0878_ _0954_ _0962_ _0963_ _1051_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_98_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6117_ _1540_ _1505_ _1575_ _2732_ _2733_ _2734_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XTAP_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_7097_ _3495_ _0283_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_432 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5247__A2 _1911_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_977 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6444__B2 _2831_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3006 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6048_ _2560_ _2664_ _2665_ _2666_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_100_465 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3017 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3028 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_160_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3039 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2305 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2316 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2327 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2338 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7244__I0 _3539_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2349 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1604 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1615 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1626 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_7999_ _0208_ net1 mod.Data_Mem.F_M.MRAM\[13\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_82_894 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_148_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7795__I1 mod.Data_Mem.F_M.MRAM\[798\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1637 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1648 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1659 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_169_46 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_1216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_167_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8536__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3981__A2 mod.Arithmetic.CN.I_in\[48\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_155_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5183__A1 _1844_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7046__S _3469_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_68_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_21 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_150_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_111_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5486__A2 _2075_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6435__A1 _2417_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_76_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8066__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7235__I0 _3531_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6038__I1 mod.Data_Mem.F_M.MRAM\[771\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2850 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_574 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2861 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_127_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2872 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_127_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4932__I _1600_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2883 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_32_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4749__A1 _0623_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2894 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_159_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6352__C _1725_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3972__A2 _0648_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7903__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_145_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5763__I _2101_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_1212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5350_ mod.Data_Mem.F_M.MRAM\[787\]\[6\] _2013_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_142_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4301_ _0901_ _0970_ _0974_ _0975_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_126_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5281_ mod.Data_Mem.F_M.MRAM\[785\]\[5\] mod.Data_Mem.F_M.MRAM\[784\]\[5\] _1942_
+ _1945_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__6123__B1 _1520_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7020_ _3242_ _3452_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4232_ _0904_ _0905_ _0906_ _0907_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_96_931 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_730 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4163_ _0658_ _0838_ _0839_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__8409__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6426__A1 _2301_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4094_ _0747_ _0765_ _0769_ _0770_ _0771_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_95_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7922_ _0148_ net1 mod.Data_Mem.F_M.MRAM\[0\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_55_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7853_ mod.Data_Mem.F_M.MRAM\[9\]\[5\] _3929_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_82_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6543__B _3107_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8559__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6804_ mod.Data_Mem.F_M.MRAM\[799\]\[6\] _3319_ _3313_ _3320_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_24_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_51_533 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_7784_ _3293_ mod.Data_Mem.F_M.MRAM\[798\]\[0\] _3889_ _3890_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4996_ _1663_ _1664_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_149_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6735_ _3269_ _3270_ _3272_ _3273_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_23_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3947_ _0624_ _0625_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_20_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_165_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6666_ _3223_ _0124_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_31_290 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8405_ _0501_ net1 mod.Data_Mem.F_M.MRAM\[787\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5617_ _1737_ _2250_ _2251_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__5165__A1 _1608_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6597_ mod.Data_Mem.F_M.MRAM\[11\]\[2\] _3189_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6901__A2 _3371_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8336_ _0432_ net1 mod.Data_Mem.F_M.MRAM\[778\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5548_ _2187_ _2188_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5960__I0 mod.Data_Mem.F_M.MRAM\[16\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_117_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6114__B1 _1809_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8267_ _0363_ net1 mod.Data_Mem.F_M.MRAM\[768\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5479_ _0025_ _2124_ _2125_ _2095_ _2126_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_105_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7218_ _3533_ mod.Data_Mem.F_M.MRAM\[2\]\[4\] _3567_ _3568_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_132_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_120_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8198_ _0083_ net2 net1 mod.I_addr\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_8_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_154_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_59_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7149_ _3526_ _0304_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_63_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4140__A2 mod.Arithmetic.CN.I_in\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8089__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6437__C _3026_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_817 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_986 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_284 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2102 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2113 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2124 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2135 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5640__A2 _2263_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_319 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1401 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2146 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2157 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1412 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2168 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1423 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2179 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1434 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_64_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4752__I _0623_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1445 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_154_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_1456 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7926__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1467 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_717 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1478 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1489 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_1160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_22_290 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3954__A2 _0630_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5583__I _1549_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5251__S1 _1915_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_97_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_739 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_145_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_78_997 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_1197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_92_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_617 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7759__I1 mod.Data_Mem.F_M.MRAM\[796\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5758__I _1588_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2680 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4850_ _1518_ _1519_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_72_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2691 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6082__C _2698_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4781_ _1174_ _1448_ _1449_ _1450_ _1451_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XTAP_1990 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6520_ _3106_ mod.Data_Mem.F_M.MRAM\[781\]\[5\] _3124_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_147_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_119_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6451_ _2258_ mod.Data_Mem.F_M.MRAM\[769\]\[2\] _3058_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_101_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_9_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5402_ _2062_ _2063_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6382_ _2895_ _2990_ _2991_ _2898_ _1866_ _2992_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_86_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_114_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8121_ mod.Data_Mem.F_M.out_data\[31\] net2 net1 mod.Arithmetic.CN.I_in\[31\] vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_114_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5333_ mod.Data_Mem.F_M.MRAM\[19\]\[6\] mod.Data_Mem.F_M.MRAM\[18\]\[6\] _1892_ _1996_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_47_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8231__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_1037 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8052_ _0261_ net1 mod.Data_Mem.F_M.MRAM\[1\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5264_ _1900_ _1928_ _1929_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_69_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7003_ _3399_ mod.Data_Mem.F_M.MRAM\[17\]\[4\] _3440_ _3441_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4215_ _0830_ _0834_ _0890_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_68_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5195_ _1621_ _1839_ _1860_ _1490_ _1861_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_84_901 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_986 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4146_ _0652_ _0657_ _0822_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_95_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8381__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4077_ _0707_ _0754_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_83_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7949__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5622__A2 _2252_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4425__A3 _0897_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7905_ _0131_ net1 mod.Data_Mem.F_M.MRAM\[28\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_43_319 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_1111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_1144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_169_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_7836_ _3907_ mod.I_addr\[2\] _3919_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_169_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_51_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_588 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4189__A2 _0851_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5386__A1 _1700_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4979_ _1646_ _1647_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_7767_ _3303_ mod.Data_Mem.F_M.MRAM\[797\]\[1\] _3878_ _3880_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_6718_ _3262_ _0137_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_7698_ mod.Data_Mem.F_M.MRAM\[793\]\[1\] _3843_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6649_ mod.Data_Mem.F_M.MRAM\[25\]\[4\] _3215_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_109_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_164_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5689__A2 _2137_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8319_ _0415_ net1 mod.Data_Mem.F_M.MRAM\[775\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_65_1104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_3_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7324__S _3625_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_717 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_160_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_115_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_59_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5779__S _1791_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_74_433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_904 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_1211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5578__I _1493_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1220 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1231 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1242 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1253 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1264 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6413__I1 mod.Data_Mem.F_M.MRAM\[1\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1275 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8104__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5377__A1 mod.Data_Mem.F_M.MRAM\[783\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1286 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_536 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1297 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_129_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_156_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__8254__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5837__C1 _2460_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_111_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4000_ mod.Arithmetic.I_out\[79\] _0677_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_66_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_66_978 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_1019 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_52_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_797 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5951_ _2162_ _2572_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_65_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4902_ _1528_ _1541_ _1571_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_80_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5882_ _2500_ _2501_ _2502_ _2503_ _2504_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_34_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7621_ _3803_ _0499_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4833_ mod.Data_Mem.F_M.src\[0\] _1502_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_61_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7552_ _3761_ _0472_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4764_ _1352_ _1361_ _1433_ _1225_ _1434_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_119_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4040__A1 _0710_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6540__C _2170_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4040__B2 _0716_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6503_ _3106_ mod.Data_Mem.F_M.MRAM\[769\]\[4\] _3107_ _3108_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_53_1085 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7483_ _3717_ _0447_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4695_ mod.Arithmetic.CN.I_in\[62\] _1366_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_146_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7208__I _3561_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6434_ _2343_ mod.Data_Mem.F_M.MRAM\[12\]\[1\] _3042_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_88_1137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_162_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6365_ _2876_ _2024_ _2715_ _2975_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_115_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5951__I _2162_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8104_ mod.Data_Mem.F_M.out_data\[14\] net2 net1 mod.Arithmetic.CN.I_in\[14\] vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_161_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5316_ mod.Data_Mem.F_M.MRAM\[19\]\[5\] mod.Data_Mem.F_M.MRAM\[18\]\[5\] _1681_ _1980_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_142_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6296_ _2144_ mod.Data_Mem.F_M.MRAM\[783\]\[4\] mod.Data_Mem.F_M.MRAM\[782\]\[4\]
+ _2267_ _2909_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_102_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_114_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_8035_ _0244_ net1 mod.Data_Mem.F_M.MRAM\[17\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__6096__A2 _1541_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7293__A1 _3612_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6983__S _3428_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5247_ _1552_ _1911_ _1884_ _1912_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_60_1001 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_1192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5843__A2 _1787_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_60_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5178_ _1526_ _1844_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_84_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4129_ _0804_ _0805_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_56_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_43_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_147_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8127__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5398__I _1522_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_169_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_24_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_325 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_7819_ mod.I_addr\[0\] mod.I_addr\[2\] mod.I_addr\[1\] _3909_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_51_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6020__A2 _2148_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8277__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_878 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_1163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_165_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_125_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_3_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4334__A2 mod.Arithmetic.CN.I_in\[67\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5531__A1 _2170_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5531__B2 _2171_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7054__S _3469_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_1092 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_503 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_161_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_1035 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_156_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_43_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4637__A3 _1062_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_904 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_606 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1050 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1061 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1072 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1083 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7229__S _3574_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1094 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6011__A2 _2618_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4940__I _1509_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4022__A1 _0696_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5770__A1 _1595_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5972__S _2528_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_939 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_7_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4480_ _1042_ _1150_ _1151_ _1152_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_128_287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6867__I mod.Data_Mem.F_M.MRAM\[6\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5373__I1 mod.Data_Mem.F_M.MRAM\[16\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5522__A1 _2161_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5522__B2 _2162_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5771__I _2395_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6150_ _1742_ _1648_ _2766_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_801 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_1007 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_823 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_83_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5101_ _1764_ _1767_ _1768_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_140_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6081_ _1756_ _2698_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_856 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_867 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_878 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5032_ _1562_ _1700_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_111_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5720__B _2280_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6535__C _3137_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6983_ _3399_ mod.Data_Mem.F_M.MRAM\[16\]\[4\] _3428_ _3429_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_81_745 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6250__A2 _1627_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5934_ _2379_ _2545_ _2554_ _2555_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_81_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_1178 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4800__A3 _1469_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5865_ _2449_ _2485_ _2486_ _2367_ _2487_ _2454_ _2488_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_21_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6538__B1 _2631_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6551__B _2103_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5946__I _2283_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4850__I _1518_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6002__A2 mod.Data_Mem.F_M.MRAM\[783\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7604_ _3793_ _0492_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__7050__I1 mod.Data_Mem.F_M.MRAM\[1\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4816_ _1395_ _1392_ _1484_ _1486_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_8584_ _0600_ net1 mod.Data_Mem.F_M.MRAM\[9\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_22_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_21_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5796_ _2417_ _1682_ _2419_ _2420_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__5167__B _1531_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6978__S _3423_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5761__A1 _1954_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4747_ _1373_ mod.Arithmetic.CN.I_in\[70\] _1416_ _1417_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_7535_ _3750_ _0466_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_108_917 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7990__RN net2 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7466_ _3603_ mod.Data_Mem.F_M.MRAM\[780\]\[0\] _3707_ _3708_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4678_ _1236_ _1255_ _1348_ _1349_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_119_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6417_ _2092_ _3026_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5513__A1 _1715_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7397_ mod.Data_Mem.F_M.MRAM\[774\]\[7\] _3672_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5364__I1 mod.Data_Mem.F_M.MRAM\[2\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5614__C _2248_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6348_ _2955_ _2956_ _2957_ _2958_ _2959_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_153_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_611 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6279_ _2891_ _1907_ _2892_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_88_355 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6474__C1 _2529_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8018_ _0227_ net1 mod.Data_Mem.F_M.MRAM\[15\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_103_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4875__I0 mod.Data_Mem.F_M.MRAM\[6\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_57_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_100 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_72_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_122 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_642 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_155 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__7041__I1 mod.Data_Mem.F_M.MRAM\[1\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_166 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_355 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_177 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_36_1080 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__4555__A2 mod.Arithmetic.CN.I_in\[58\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5752__A1 _2106_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_158_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_126_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5504__A1 _1791_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4307__A2 _0829_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6687__I _3239_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5591__I _1606_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_137_82 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_1207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_1040 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_153_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6480__A2 _3085_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8442__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4491__A1 _1075_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_35_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_745 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4871__S _1514_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_907 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3980_ _0655_ _0656_ _0657_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XPHY_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_22_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_16_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_62_288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5991__A1 _2414_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8592__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5650_ _2281_ mod.Data_Mem.F_M.MRAM\[29\]\[1\] _2282_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_15_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4601_ _1149_ _1270_ _1271_ _1272_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_129_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4546__A2 _1212_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5581_ _2213_ _2179_ _2215_ _2218_ _2219_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_129_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7320_ _3615_ mod.Data_Mem.F_M.MRAM\[770\]\[4\] _3623_ _3630_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4532_ _1101_ _1204_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_8_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_50_1088 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7251_ _3587_ _0345_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4463_ _0642_ mod.Arithmetic.CN.I_in\[60\] _1136_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6202_ _2681_ _2813_ _2816_ _2817_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_125_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7182_ _3546_ _0317_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4394_ _1058_ _1060_ _1065_ _1066_ _1067_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
XFILLER_131_249 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6133_ _2682_ _2747_ _2748_ _2084_ _2749_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XTAP_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_642 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_675 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6064_ _1840_ _2402_ _1535_ _2681_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_86_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_61_1151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5015_ _1681_ _1682_ _1683_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__6038__S _2339_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4482__A1 _0988_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_1195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2509 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6223__A2 _2685_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1808 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1819 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6966_ _3403_ mod.Data_Mem.F_M.MRAM\[15\]\[6\] _3414_ _3418_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_54_789 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4234__A1 _0619_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5917_ _2506_ mod.Data_Mem.F_M.MRAM\[788\]\[4\] _2537_ _2538_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_22_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6897_ _3334_ _3371_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_22_642 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_50_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5848_ _2428_ _1784_ _2429_ _2470_ _2471_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__5034__I0 mod.Data_Mem.F_M.MRAM\[773\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4537__A2 mod.Arithmetic.CN.I_in\[44\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8567_ _0071_ net1 mod.Data_Mem.F_M.out_data\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5779_ mod.Data_Mem.F_M.MRAM\[784\]\[0\] mod.Data_Mem.F_M.MRAM\[785\]\[0\] _1791_
+ _2404_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_166_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_120_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7518_ _3725_ mod.Data_Mem.F_M.MRAM\[782\]\[4\] _3739_ _3740_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_108_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_8498_ _0002_ net1 mod.Data_Mem.F_M.out_data\[74\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__8315__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_107_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7449_ mod.Data_Mem.F_M.MRAM\[778\]\[1\] _3698_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_107_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_162_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_964 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8465__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_49_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6447__C1 _2469_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6837__I1 mod.Data_Mem.F_M.MRAM\[769\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8140__RN net2 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_91_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_29_252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6175__C _2743_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4863__I3 _1520_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6214__A2 _2828_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4776__A2 _1321_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5973__A1 _2510_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5973__B2 _2565_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_8_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_158_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5725__A1 _2068_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4528__A2 _1140_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5725__B2 _2168_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_500 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5328__I1 _1988_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_154_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6150__A1 _1742_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_1151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_1184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7242__S _3579_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_1059 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8131__RN net2 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_678 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4464__A1 _0923_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_82_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6205__A2 _1772_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6820_ mod.Data_Mem.F_M.MRAM\[789\]\[5\] _3329_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_51_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7982__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_726 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6751_ _3282_ _0150_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5964__A1 _2558_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3963_ _0613_ _0640_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_50_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7005__I1 mod.Data_Mem.F_M.MRAM\[17\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_1144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5702_ _2203_ mod.Data_Mem.F_M.MRAM\[797\]\[5\] _2330_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_6682_ _3230_ _3232_ _3235_ _3236_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_52_1117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_1188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8338__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8198__RN net2 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8421_ _0517_ net1 mod.Data_Mem.F_M.MRAM\[790\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5633_ _1875_ _2266_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_148_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6321__S _2044_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5564_ _2096_ _2203_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_8352_ _0448_ net1 mod.Data_Mem.F_M.MRAM\[781\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_7303_ _3618_ mod.Data_Mem.F_M.MRAM\[768\]\[6\] _3608_ _3619_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4515_ _1166_ _1184_ _1186_ _1187_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
X_8283_ _0379_ net1 mod.Data_Mem.F_M.MRAM\[771\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5495_ _2138_ mod.Data_Mem.F_M.MRAM\[798\]\[4\] _2139_ _2140_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XANTENNA__8488__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_588 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7234_ _3577_ _0338_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4446_ _0828_ _0930_ _0928_ _1114_ _1119_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
XANTENNA__6141__A1 _2192_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7165_ _3255_ _3537_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_160_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4377_ _0962_ _0963_ _0877_ _0954_ _1050_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_101_901 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_113_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_112_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6116_ _2714_ _2733_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_98_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7096_ mod.Data_Mem.F_M.MRAM\[23\]\[3\] _3495_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_112_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_461 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6047_ _2214_ mod.Data_Mem.F_M.MRAM\[20\]\[7\] _2665_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_74_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8122__RN net2 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6444__A2 _3048_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3007 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3018 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4455__A1 _0640_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_3029 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2306 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_54_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2317 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2328 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2339 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6790__I _3308_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7244__I1 mod.Data_Mem.F_M.MRAM\[30\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1605 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4207__A1 _0813_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1616 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_7998_ mod.P2.dest_reg1\[8\] net2 net1 mod.P2.dest_reg\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_42_726 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1627 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1638 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1649 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5955__A1 _2410_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4758__A2 _1427_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6949_ _3295_ _3407_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_41_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_169_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_781 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7835__B _3916_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_154_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_167_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_108_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5183__A2 _1848_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_136_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_68_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_897 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_1168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6132__A1 _2183_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_33 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_155_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_111_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4694__A1 _1249_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5318__S0 _1527_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8113__RN net2 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6435__A2 mod.Data_Mem.F_M.MRAM\[13\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_83 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_64_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4446__A1 _0828_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_1220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7235__I1 mod.Data_Mem.F_M.MRAM\[30\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_166_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6199__A1 _2425_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2840 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2851 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6199__B2 _2448_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5246__I0 _1904_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5310__S _1968_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2862 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2873 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2884 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4749__A2 mod.Arithmetic.CN.I_in\[70\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2895 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6994__I0 _3386_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_159_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6746__I0 _3249_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_160_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4300_ _0972_ _0973_ _0974_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_5280_ _1941_ _1943_ _1944_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__6123__A1 _1795_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6123__B2 _1713_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4231_ _0837_ _0848_ _0906_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_102_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_49_1090 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5882__B1 _2502_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4162_ _0635_ mod.Arithmetic.CN.I_in\[49\] _0838_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_96_943 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_645 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7623__A1 _3312_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8104__RN net2 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_678 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4093_ _0763_ _0764_ _0748_ _0770_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_55_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8010__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4437__A1 _0993_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7921_ _0147_ net1 mod.Data_Mem.F_M.MRAM\[0\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_55_339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7852_ _3928_ _0604_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_36_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6803_ _3318_ _3319_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__8160__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6985__I0 _3416_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7783_ _3888_ _3889_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_23_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4995_ _1525_ _1663_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_51_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6734_ _3271_ _3272_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_3946_ _0623_ _0624_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_56_1094 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_104_1004 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6665_ mod.Data_Mem.F_M.MRAM\[27\]\[4\] _3223_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6737__I0 _3228_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_1037 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8404_ _0500_ net1 mod.Data_Mem.F_M.MRAM\[787\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_149_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5616_ _1746_ mod.Data_Mem.F_M.MRAM\[31\]\[7\] mod.Data_Mem.F_M.MRAM\[30\]\[7\] _2187_
+ _2250_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_30_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5165__A2 _1830_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6596_ _3188_ _0089_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__7878__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8335_ _0431_ net1 mod.Data_Mem.F_M.MRAM\[777\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5547_ _1914_ _2187_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__5960__I1 mod.Data_Mem.F_M.MRAM\[17\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6114__A1 mod.Data_Mem.F_M.MRAM\[1\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6114__B2 mod.Data_Mem.F_M.MRAM\[0\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8266_ _0362_ net1 mod.Data_Mem.F_M.MRAM\[768\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5478_ mod.Data_Mem.F_M.MRAM\[798\]\[2\] mod.Data_Mem.F_M.MRAM\[799\]\[2\] _1890_
+ _2125_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_7217_ _3561_ _3567_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_4429_ _1095_ _1101_ _1102_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__6785__I net5 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8197_ _0082_ net2 net1 mod.I_addr\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_8_1213 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7148_ _3523_ mod.Data_Mem.F_M.MRAM\[12\]\[0\] _3525_ _3526_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_98_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4140__A3 _0709_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_150_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7079_ _3486_ _0274_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_101_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4428__A1 _1096_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_1117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_497 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2103 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8503__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2114 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2125 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2136 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5640__A3 _2272_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2147 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1402 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2158 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5228__I0 mod.Data_Mem.F_M.MRAM\[19\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1413 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1424 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2169 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1435 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6976__I0 _3393_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1446 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_159_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1468 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1479 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_147_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_80_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_161_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_1025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_155_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6353__A1 _2951_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_124_801 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_6_468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_159_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_65 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6105__A1 _2620_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6105__B2 _2162_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6695__I _3245_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__8033__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5305__S _1968_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__4419__A1 _0893_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7520__S _3739_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5616__B1 mod.Data_Mem.F_M.MRAM\[30\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_161_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8183__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4943__I _1567_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_166_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_61_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2670 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2681 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2692 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4780_ _1309_ _1317_ _1450_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_53_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1980 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1991 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_118_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6344__A1 _1635_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6450_ _2696_ mod.Data_Mem.F_M.MRAM\[780\]\[2\] _2382_ _3057_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_5401_ _2061_ _2062_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_62_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_6381_ _2051_ _2052_ _1881_ _2991_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_103_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_161_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_103_1092 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5332_ mod.Data_Mem.F_M.MRAM\[21\]\[6\] mod.Data_Mem.F_M.MRAM\[20\]\[6\] _1892_ _1995_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_8120_ mod.Data_Mem.F_M.out_data\[30\] net2 net1 mod.Arithmetic.CN.I_in\[30\] vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XANTENNA__5723__B _2217_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8051_ _0260_ net1 mod.Data_Mem.F_M.MRAM\[1\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5263_ _1902_ _1912_ _1926_ _1927_ _1629_ _1928_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_138_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5215__S _1879_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4658__A1 _1208_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4658__B2 _1217_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7002_ _3434_ _3440_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_4214_ _0836_ _0887_ _0888_ _0889_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_102_539 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5194_ _1721_ _1850_ _1859_ _1860_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_60_1216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8526__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4145_ _0621_ _0656_ _0820_ _0821_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__5607__B1 _1749_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4076_ _0750_ _0751_ _0704_ _0752_ _0753_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XANTENNA__5083__A1 mod.Data_Mem.F_M.MRAM\[22\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7904_ _0130_ net1 mod.Data_Mem.F_M.MRAM\[28\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_93_1014 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7835_ _3175_ _3918_ _3916_ _0598_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_58_1156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_1058 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5386__A2 _2047_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7766_ _3879_ _0568_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4978_ _1593_ _1646_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6717_ mod.Data_Mem.F_M.MRAM\[10\]\[1\] _3262_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5684__I _1691_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_165_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_7697_ _3842_ _0536_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_137_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6648_ _3214_ _0115_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6335__A1 _1635_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_166_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_153_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_124_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6579_ _3177_ _0083_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__8056__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7605__S _3787_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8318_ _0414_ net1 mod.Data_Mem.F_M.MRAM\[775\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_105_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_8249_ _0345_ net1 mod.Data_Mem.F_M.MRAM\[31\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_133_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_78_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_604 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_968 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6464__B _2073_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_607 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1210 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_43_843 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1232 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1243 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_651 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1254 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1265 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_91_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1276 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5377__A2 _1673_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1287 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1298 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6326__A1 mod.Data_Mem.F_M.MRAM\[13\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6326__B2 mod.Data_Mem.F_M.MRAM\[12\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7515__S _3734_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4003__I mod.Arithmetic.CN.I_in\[19\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_1216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8549__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4938__I _1606_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5035__S _1692_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5837__C2 _2170_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_78_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7250__S _3585_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5065__A1 _1730_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5950_ _2266_ mod.Data_Mem.F_M.MRAM\[4\]\[4\] _2571_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_34_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3190 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_80_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4901_ _1566_ _1569_ _1570_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5881_ _2376_ _2503_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_7620_ _3765_ mod.Data_Mem.F_M.MRAM\[787\]\[3\] _3801_ _3803_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__7601__I1 mod.Data_Mem.F_M.MRAM\[786\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4832_ _1500_ _1501_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6565__A1 _3017_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5368__A2 _2029_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7551_ _3718_ mod.Data_Mem.F_M.MRAM\[784\]\[0\] _3760_ _3761_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_18_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_53_1053 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4763_ _1251_ _1354_ mod.Arithmetic.CN.I_in\[54\] _1433_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_147_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_144_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8079__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6502_ _2102_ _3107_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6317__A1 _2718_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7482_ _3620_ mod.Data_Mem.F_M.MRAM\[780\]\[7\] _3713_ _3717_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4694_ _1249_ _1253_ _1364_ _1365_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_107_609 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_1127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6433_ _2626_ _3032_ _3040_ _3041_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_106_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5009__I _1676_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7117__I0 _3456_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6364_ _1585_ _2026_ _2974_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_8103_ mod.Data_Mem.F_M.out_data\[13\] net2 net1 mod.Arithmetic.CN.I_in\[13\] vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_5315_ mod.Data_Mem.F_M.MRAM\[21\]\[5\] mod.Data_Mem.F_M.MRAM\[20\]\[5\] _1968_ _1979_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_6295_ mod.Data_Mem.F_M.MRAM\[13\]\[4\] _2901_ _2902_ mod.Data_Mem.F_M.MRAM\[12\]\[4\]
+ _2907_ _2908_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_0_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7916__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8034_ _0243_ net1 mod.Data_Mem.F_M.MRAM\[17\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__7293__A2 _3606_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5246_ _1904_ _1905_ _1907_ _1909_ _1910_ _1805_ _1911_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_102_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_1013 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_615 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5177_ _1745_ _1842_ _1843_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_56_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_69_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4128_ _0803_ _0804_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_44_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4059_ _0735_ _0730_ _0736_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__4803__A1 _1444_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_71_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_80_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_52_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_326 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_7818_ mod.I_addr\[4\] mod.I_addr\[6\] mod.I_addr\[5\] mod.I_addr\[7\] _3908_ vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_52_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__6556__A1 _3021_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7749_ _3869_ _0561_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_123_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_1175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6308__A1 _2869_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7108__I0 _3445_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_152_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_642 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_1082 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_3_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6973__I _3422_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_946 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5589__I _1549_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5598__A2 mod.Data_Mem.F_M.MRAM\[799\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1040 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_35_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1051 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_1075 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8221__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1062 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_71_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1073 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1084 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_163_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_129_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7309__I _3622_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_156_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7347__I0 _3618_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_907 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_11_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5770__A2 _1554_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8371__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7939__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5522__A2 mod.Data_Mem.F_M.MRAM\[30\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_1182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_1084 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_48_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5100_ _1707_ mod.Data_Mem.F_M.MRAM\[771\]\[2\] _1766_ _1767_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_97_323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_1019 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6080_ _2696_ mod.Data_Mem.F_M.MRAM\[14\]\[0\] mod.Data_Mem.F_M.MRAM\[15\]\[0\] _2517_
+ _2697_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_846 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_868 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5031_ _1672_ _1699_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_100_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_879 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_25_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_81_724 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6982_ _3422_ _3428_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_65_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5933_ _2434_ _2553_ _2554_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_1157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_1104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_1153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_80_278 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_1126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5864_ mod.Data_Mem.F_M.MRAM\[18\]\[2\] mod.Data_Mem.F_M.MRAM\[19\]\[2\] _2452_ _2487_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_34_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6538__A1 _2447_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_1017 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6538__B2 _2642_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7603_ _3778_ mod.Data_Mem.F_M.MRAM\[786\]\[4\] _3787_ _3793_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4815_ _1395_ _1392_ _1484_ _1485_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
X_8583_ _0599_ net1 mod.Instr_Mem.instruction\[23\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5795_ _2418_ mod.Data_Mem.F_M.MRAM\[787\]\[1\] _2419_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_7534_ _3749_ mod.Data_Mem.F_M.MRAM\[783\]\[2\] _3745_ _3750_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4746_ mod.Arithmetic.CN.I_in\[69\] _1376_ _1416_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_7465_ _3706_ _3707_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_107_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4677_ _1237_ _1254_ _1348_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_107_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_162_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6416_ _3014_ _3019_ _3024_ _3025_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__5513__A2 mod.Data_Mem.F_M.MRAM\[799\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_1200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7396_ _3671_ _0406_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_89_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6994__S _3435_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4578__I mod.Arithmetic.CN.I_in\[61\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6347_ _2012_ _1988_ _2739_ _2958_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_131_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6278_ _2228_ _2891_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_131_987 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6474__B1 _3006_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_678 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8017_ _0226_ net1 mod.Data_Mem.F_M.MRAM\[15\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__6793__I net7 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6474__C2 _2510_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5229_ _1813_ _1894_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_88_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5029__A1 _1674_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8244__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6777__A1 _3294_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_426 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4252__A2 _0921_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_71_278 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_112 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_53_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6529__A1 _2534_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_123 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_24_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_134 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_80_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_145 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_169_166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8394__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_167 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_169_177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5201__A1 _1757_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_178 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_189 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__5201__B2 _1721_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4555__A3 mod.Arithmetic.CN.I_in\[59\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5752__A2 _2376_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_165_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5504__A2 mod.Data_Mem.F_M.MRAM\[31\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_153_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_761 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_94_348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_787 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4491__A2 _1076_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5112__I _1579_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_3 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_44_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5440__A1 _2072_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_971 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_278 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_50_429 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4600_ _1152_ _1259_ _1271_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__4546__A3 _1217_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5580_ _2061_ mod.Data_Mem.F_M.MRAM\[30\]\[3\] _2217_ _2218_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_157_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_117_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4531_ _1202_ _1203_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_144_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_7250_ _1632_ _3303_ _3585_ _3587_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4462_ _0635_ _1017_ _1134_ _1135_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_116_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8117__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6201_ _1661_ _2814_ _2815_ _2775_ _2816_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_104_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4393_ _0642_ _0959_ _1062_ _1055_ _1066_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
X_7181_ mod.Data_Mem.F_M.MRAM\[22\]\[5\] _3546_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_98_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_610 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6132_ _2183_ _2689_ _2748_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_140_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_643 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5259__A1 _1834_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_998 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_615 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6063_ _2534_ _2662_ _2680_ _2414_ _0063_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8267__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_1163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5014_ mod.Data_Mem.F_M.MRAM\[786\]\[1\] _1682_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__6059__I0 mod.Data_Mem.F_M.MRAM\[14\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5022__I _1522_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1809 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6965_ _3417_ _0229_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4234__A2 _0661_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4861__I _1529_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5916_ _2428_ mod.Data_Mem.F_M.MRAM\[789\]\[4\] _2537_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_35_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6896_ _3370_ _0207_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__3993__A1 _0652_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6989__S _3428_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5847_ _2358_ mod.Data_Mem.F_M.MRAM\[789\]\[2\] _2470_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_146_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_985 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5034__I1 mod.Data_Mem.F_M.MRAM\[772\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8566_ _0070_ net1 mod.Data_Mem.F_M.out_data\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5778_ _2402_ _2403_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_120_1213 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_147_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7517_ _3733_ _3739_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_4729_ _1279_ _1397_ _1398_ _1399_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_8497_ _0001_ net1 mod.Data_Mem.F_M.out_data\[73\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_163_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_7448_ _3697_ _0432_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_135_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5498__A1 _1778_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7379_ mod.Data_Mem.F_M.MRAM\[773\]\[6\] _3663_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__7613__S _3798_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4101__I _0746_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7840__C _3916_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6447__B1 _3006_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6447__C2 _3023_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_464 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3940__I _0617_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5670__A1 _2270_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_584 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_60_716 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_73_1001 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_610 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5973__A2 _2591_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6191__C _2763_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_125_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_985 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6922__A1 mod.Data_Mem.F_M.dest\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5725__A2 _2347_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6698__I net7 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_126_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5328__I2 _1989_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6150__A2 _1648_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4161__A1 _0660_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_1163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_1196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_1049 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_819 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4464__A2 _1019_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_169_1073 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_36_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_35_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6750_ _3256_ mod.Data_Mem.F_M.MRAM\[0\]\[6\] _3279_ _3282_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_17_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3962_ _0637_ mod.Arithmetic.CN.I_in\[24\] _0638_ _0639_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XANTENNA_output9_I net9 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5964__A2 _2580_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3975__A1 _0651_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5701_ _2325_ _2327_ _2328_ _2329_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_92_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_91_1156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6681_ _3234_ _3235_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_8420_ _0516_ net1 mod.Data_Mem.F_M.MRAM\[790\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5632_ _2264_ mod.Data_Mem.F_M.MRAM\[29\]\[0\] _2265_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_8351_ _0447_ net1 mod.Data_Mem.F_M.MRAM\[780\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5563_ _2201_ _2202_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_7302_ _3318_ _3618_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_145_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4514_ _1185_ _1093_ _1186_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_8282_ _0378_ net1 mod.Data_Mem.F_M.MRAM\[771\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5494_ _1677_ mod.Data_Mem.F_M.MRAM\[799\]\[4\] _2139_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_117_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8511__187 net187 vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
X_7233_ _3529_ mod.Data_Mem.F_M.MRAM\[30\]\[2\] _3574_ _3577_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4445_ _1112_ _1117_ _1118_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__5017__I _1518_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6141__A2 _2689_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7164_ _3536_ _0309_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_59_805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4376_ _0966_ _0965_ _1049_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__6557__B _1757_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6115_ mod.Data_Mem.F_M.MRAM\[7\]\[0\] mod.Data_Mem.F_M.MRAM\[6\]\[0\] _1707_ _2732_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4856__I _1524_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_7095_ _3494_ _0282_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_462 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_473 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6046_ _2620_ mod.Data_Mem.F_M.MRAM\[21\]\[7\] _2664_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_86_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3008 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3019 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5652__A1 _2283_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4455__A2 mod.Arithmetic.ACTI.x\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_893 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2307 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_148_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2318 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_66_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2329 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1606 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_7997_ mod.P2.dest_reg1\[4\] net2 net1 mod.P2.dest_reg\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XANTENNA__5687__I _2267_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4207__A2 _0715_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_1018 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1617 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_26_278 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_429 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1639 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6948_ _3406_ _0223_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5955__A2 _2570_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_248 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_169_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_169_48 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6879_ mod.Data_Mem.F_M.MRAM\[6\]\[7\] _3362_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_70_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_168_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5636__B _2268_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8549_ _0053_ net1 mod.Data_Mem.F_M.out_data\[29\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_120_1021 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_108_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8432__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5355__C _1822_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_162_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6132__A2 _2689_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4143__A1 _0802_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_462 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8582__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5891__A1 _2512_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_150_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_77_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_40 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_49_326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5318__S1 _1795_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4446__A2 _0930_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_690 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2830 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_40_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_1107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2841 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6199__A2 mod.Data_Mem.F_M.MRAM\[22\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5597__I _1811_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2852 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2863 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_32_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2874 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2885 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2896 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6994__I1 mod.Data_Mem.F_M.MRAM\[17\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7518__S _3739_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4006__I mod.Arithmetic.I_out\[74\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6746__I1 mod.Data_Mem.F_M.MRAM\[0\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_9_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_843 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_127_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4382__A1 _0844_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_154_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_99_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6123__A2 _1516_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4134__A1 _0646_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_248 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4230_ _0837_ _0848_ _0905_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_68_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5882__A1 _2500_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5882__B2 _2503_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4161_ _0660_ _0667_ _0837_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_68_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4092_ _0754_ _0766_ _0767_ _0768_ _0769_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_95_465 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4437__A2 _0999_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7920_ _0146_ net1 mod.Data_Mem.F_M.MRAM\[0\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__6891__I mod.Data_Mem.F_M.MRAM\[4\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_178 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7851_ mod.Data_Mem.F_M.MRAM\[9\]\[4\] _3928_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_63_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8305__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6802_ net9 _3318_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_1_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_7782_ _3294_ _3298_ _3446_ _3888_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__5300__I _1724_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4994_ mod.Data_Mem.F_M.MRAM\[22\]\[1\] _1661_ _1531_ _1662_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__6985__I1 mod.Data_Mem.F_M.MRAM\[16\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6733_ mod.Data_Mem.F_M.dest\[4\] mod.Data_Mem.F_M.dest\[2\] _3271_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_23_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3945_ _0622_ _0623_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__8455__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6664_ _3222_ _0123_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6737__I1 mod.Data_Mem.F_M.MRAM\[0\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8403_ _0499_ net1 mod.Data_Mem.F_M.MRAM\[787\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5615_ _2225_ _2246_ _2249_ _2177_ _0046_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
X_6595_ mod.Data_Mem.F_M.MRAM\[11\]\[1\] _3188_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6362__A2 _2964_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8334_ _0430_ net1 mod.Data_Mem.F_M.MRAM\[777\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_118_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5546_ _1602_ _2186_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_117_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_8265_ _0361_ net1 mod.Data_Mem.F_M.MRAM\[768\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_144_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5477_ mod.Data_Mem.F_M.MRAM\[30\]\[2\] mod.Data_Mem.F_M.MRAM\[31\]\[2\] _1510_ _2124_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__6114__A2 _1539_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7163__S _3534_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7216_ _3566_ _0331_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4428_ _1096_ _1100_ _1101_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_8196_ _0081_ net2 net1 mod.I_addr\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_160_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_99_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7147_ _3524_ _3525_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_48_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4359_ _0781_ _0799_ _1032_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_98_270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7078_ mod.Data_Mem.F_M.MRAM\[21\]\[2\] _3486_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_59_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6029_ _2630_ _2647_ _0062_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_39_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2104 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2115 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2126 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2137 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2148 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5228__I1 mod.Data_Mem.F_M.MRAM\[18\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1403 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2159 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1414 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_64_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4027__S _0703_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1425 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1436 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5210__I _1646_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1447 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6050__A1 _2129_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1458 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1469 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_1184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_167_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_13_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_10_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_843 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_108_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_124_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_163_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7972__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5164__I0 mod.Data_Mem.F_M.MRAM\[787\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_1155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_1177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8328__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5616__A1 _1746_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4419__A2 _0980_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8098__RN net2 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5616__B2 _2187_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_690 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_969 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_79_1051 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2660 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2671 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8478__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2682 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6041__A1 _2548_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2693 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_21_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1970 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1981 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1992 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7248__S _3585_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_159_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6344__A2 _1990_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5400_ _2060_ _2061_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_103_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6380_ mod.Data_Mem.F_M.MRAM\[789\]\[7\] mod.Data_Mem.F_M.MRAM\[791\]\[7\] mod.Data_Mem.F_M.MRAM\[790\]\[7\]
+ mod.Data_Mem.F_M.MRAM\[788\]\[7\] _1915_ _2383_ _2990_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__5552__B1 _1809_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_155_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5331_ mod.Data_Mem.F_M.MRAM\[23\]\[6\] mod.Data_Mem.F_M.MRAM\[22\]\[6\] _1708_ _1994_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_126_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_1055 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4107__A1 _0730_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8050_ _0259_ net1 mod.Data_Mem.F_M.MRAM\[1\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_47_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5262_ _1653_ _1927_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_69_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_69_911 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7001_ _3439_ _0243_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_69_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4213_ _0825_ _0849_ _0888_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_102_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5193_ _1642_ _1854_ _1858_ _1859_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_68_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4144_ mod.Arithmetic.CN.I_in\[32\] _0820_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_95_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8089__RN net2 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5607__B2 mod.Data_Mem.F_M.MRAM\[796\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4075_ _0630_ _0752_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__5083__A2 _1749_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6280__A1 _2718_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_7903_ _0129_ net1 mod.Data_Mem.F_M.MRAM\[28\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_58_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_822 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7834_ _0080_ _3171_ _3918_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__6958__I1 mod.Data_Mem.F_M.MRAM\[15\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_1168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_7765_ _3293_ mod.Data_Mem.F_M.MRAM\[797\]\[0\] _3878_ _3879_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4977_ _1644_ _1645_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6716_ _3261_ _0136_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4594__A1 _1031_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7696_ mod.Data_Mem.F_M.MRAM\[793\]\[0\] _3842_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5218__S0 _1881_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_149_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6647_ mod.Data_Mem.F_M.MRAM\[25\]\[3\] _3214_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4346__A1 _0813_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7995__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5543__B1 _1640_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_146_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6578_ _3175_ _3176_ _3177_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_69_1220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8317_ _0413_ net1 mod.Data_Mem.F_M.MRAM\[775\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_105_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5529_ _1915_ _2170_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_3_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_145_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6099__A1 _2195_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_1128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8248_ _0344_ net1 mod.Data_Mem.F_M.MRAM\[31\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_78_207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_161_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_121_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5846__A1 _2424_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8179_ _0289_ net1 mod.Data_Mem.F_M.MRAM\[3\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_19_307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7599__A1 _3612_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_936 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_284 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1200 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4980__S _1647_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1211 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1222 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6559__C1 _2650_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1233 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1255 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1266 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6480__B _3047_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1288 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1299 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5808__C _2431_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_155_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8000__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4337__A1 _0641_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_610 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5316__S _1681_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5543__C _2182_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7826__A2 _3911_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5837__A1 _2458_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8150__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5837__B2 _2459_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5115__I _1518_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_730 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7531__S _3745_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_860 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7330__I _3635_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_755 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5065__A2 _1731_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6262__A1 _1655_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7868__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5986__S _1686_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3180 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4900_ mod.Data_Mem.F_M.MRAM\[773\]\[0\] mod.Data_Mem.F_M.MRAM\[772\]\[0\] _1568_
+ _1569_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_3191 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5880_ mod.Data_Mem.F_M.MRAM\[784\]\[3\] mod.Data_Mem.F_M.MRAM\[785\]\[3\] _2339_
+ _2502_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_61_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6014__A1 _2512_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2490 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4831_ mod.Data_Mem.F_M.src\[2\] _1500_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_60_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_1010 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_1021 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7550_ _3759_ _3760_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_4762_ _1410_ _1429_ _1431_ _1432_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_105_1133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6501_ _2203_ _3106_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_140_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7481_ _3716_ _0446_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4693_ _1240_ _1248_ _1364_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_101_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6432_ _1965_ _3039_ _3040_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_128_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_161_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_115_610 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6363_ _2866_ _2973_ _0070_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__7117__I1 mod.Data_Mem.F_M.MRAM\[3\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5226__S _1890_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8102_ mod.Data_Mem.F_M.out_data\[12\] net2 net1 mod.Arithmetic.CN.I_in\[12\] vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_5314_ mod.Data_Mem.F_M.MRAM\[23\]\[5\] mod.Data_Mem.F_M.MRAM\[22\]\[5\] _1568_ _1978_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_6294_ _2903_ _2906_ _2907_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_130_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_88_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8033_ _0242_ net1 mod.Data_Mem.F_M.MRAM\[17\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5245_ _1644_ _1910_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_69_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5176_ _1840_ mod.Data_Mem.F_M.MRAM\[775\]\[3\] _1841_ _1842_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_84_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_1036 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4127_ _0633_ mod.Arithmetic.CN.I_in\[17\] _0803_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_84_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_969 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4058_ _0731_ _0735_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_71_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_43_129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_149_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6005__A1 _2062_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_327 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_7817_ mod.I_addr\[3\] _3907_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XPHY_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__6800__I0 mod.Data_Mem.F_M.MRAM\[799\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_1110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8023__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7748_ _3747_ mod.Data_Mem.F_M.MRAM\[796\]\[1\] _3867_ _3869_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_137_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7679_ _3833_ _0527_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_71_1187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4104__I mod.Arithmetic.ACTI.x\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4319__A1 _0929_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_153_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5367__I0 _2024_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8173__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5644__B _2268_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3943__I _0620_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7108__I1 mod.Data_Mem.F_M.MRAM\[3\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_156_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_79_505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5819__A1 _2440_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_85 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_1059 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6492__A1 _2511_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7150__I _3239_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_714 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_90_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_43_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1030 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1052 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_674 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1085 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1096 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_169_893 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_50_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__8516__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_168_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7347__I1 mod.Data_Mem.F_M.MRAM\[771\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4014__I mod.Arithmetic.CN.I_in\[20\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_167_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_156_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_429 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6180__B1 _2202_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_1194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_1096 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_836 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7261__S _3590_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_858 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5030_ mod.Data_Mem.F_M.MRAM\[799\]\[1\] _1673_ _1697_ _1698_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_97_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_914 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_711 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_66_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6235__A1 _2160_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6981_ _3427_ _0235_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_20_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4097__I0 mod.Arithmetic.CN.I_in\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_939 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6330__S1 _2759_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_682 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8046__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5932_ _2423_ _2546_ _2547_ _2464_ _2552_ _2553_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_34_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5863_ mod.Data_Mem.F_M.MRAM\[2\]\[2\] mod.Data_Mem.F_M.MRAM\[3\]\[2\] _1954_ _2486_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__6538__A2 _2337_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7602_ _3792_ _0491_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_61_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4814_ _1396_ _1483_ _1484_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__4549__A1 _1122_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5746__B1 _2365_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8582_ _0598_ net1 mod.Instr_Mem.instruction\[22\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5794_ _1517_ _2418_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_166_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8196__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7533_ _3305_ _3749_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_119_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4745_ _0622_ mod.Arithmetic.CN.I_in\[71\] _1415_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_7464_ _3269_ _3705_ _3374_ _3706_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_119_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4676_ _1346_ _1347_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_134_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6415_ _3021_ _2359_ _3022_ _3023_ _3009_ _2368_ _3024_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_1
X_7395_ mod.Data_Mem.F_M.MRAM\[774\]\[6\] _3671_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_66_1212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6346_ _2876_ _1987_ _2957_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_102_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6277_ _1826_ _1909_ _2890_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_8016_ _0225_ net1 mod.Data_Mem.F_M.MRAM\[15\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__6474__A1 _3026_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5228_ mod.Data_Mem.F_M.MRAM\[19\]\[4\] mod.Data_Mem.F_M.MRAM\[18\]\[4\] _1892_ _1893_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_76_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6474__B2 _2523_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5159_ _1804_ _1824_ _1825_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_56_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_57_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5029__A2 _1696_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6226__A1 _1585_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_714 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_574 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6777__A2 _3296_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4788__A1 _1234_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_102 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_73_1216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_113 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__8539__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_80_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3938__I _0615_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_135 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_13_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4035__S _0702_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_146 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__5358__C _1629_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_157 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__5201__A2 mod.Data_Mem.F_M.MRAM\[15\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4555__A4 _1136_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__4960__A1 _1625_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_21_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_4_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_985 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_79_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_432 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5899__S0 _1918_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_43_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_711 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8069__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_4 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_50_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5440__A2 _2074_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_983 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4453__B _0645_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7906__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_148_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_50_1002 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_1013 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_1201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4530_ mod.Arithmetic.CN.I_in\[44\] _1202_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_89_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_1068 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_7_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4461_ mod.Arithmetic.CN.I_in\[60\] _1134_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6200_ _2761_ _1752_ _2815_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__6099__C _2715_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4703__A1 mod.Arithmetic.CN.I_in\[67\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7180_ _3545_ _0316_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4392_ _1061_ _1063_ _1064_ _0871_ _1065_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_113_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_611 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6131_ _2169_ _2745_ _2746_ _2747_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_611 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_98_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5259__A2 _1921_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6456__A1 _3003_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6062_ _2531_ _2671_ _2679_ _2680_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_100_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_677 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5013_ _1676_ _1681_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_100_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_1175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6208__A1 _2779_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6059__I1 mod.Data_Mem.F_M.MRAM\[15\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_54_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_38_287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_93_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_393 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6964_ _3416_ mod.Data_Mem.F_M.MRAM\[15\]\[5\] _3414_ _3417_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_54_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4234__A3 mod.Arithmetic.CN.I_in\[64\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5915_ _2440_ _2536_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6895_ mod.Data_Mem.F_M.MRAM\[4\]\[7\] _3370_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_107_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6134__I _2685_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3993__A2 _0657_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5846_ _2424_ _1792_ _2468_ _2469_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_167_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_1058 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5195__A1 _1621_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8565_ _0069_ net1 mod.Data_Mem.F_M.out_data\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5777_ _2008_ _1548_ _2402_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__7166__S _3534_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7516_ _3738_ _0459_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4728_ _1282_ _1387_ _1398_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__4942__A1 _1608_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8496_ _0000_ net1 mod.Data_Mem.F_M.out_data\[72\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_108_738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_162_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_7447_ mod.Data_Mem.F_M.MRAM\[778\]\[0\] _3697_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4659_ mod.Arithmetic.CN.I_in\[37\] _1330_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_123_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5498__A2 mod.Data_Mem.F_M.MRAM\[798\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7378_ _3662_ _0397_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_66_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_150_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_1042 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6329_ mod.Data_Mem.F_M.MRAM\[781\]\[5\] _2751_ _2157_ mod.Data_Mem.F_M.MRAM\[780\]\[5\]
+ _2940_ _2941_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_89_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8211__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_817 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6447__A1 _3005_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6447__B2 _2466_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_153_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_130_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_88_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5670__A2 _2127_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8361__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_213 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7929__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6472__C _3077_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_1171 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_1193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_38_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_964 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5186__A1 _1647_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_157_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6383__B1 _2989_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_154_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5328__I3 _1990_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_153_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_107_771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_79_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4161__A2 _0667_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5324__S _1873_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_79_187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5110__A1 _1759_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7238__I0 _3533_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_574 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_91_820 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_169_1052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_36_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_533 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_393 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6382__C _1866_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3961_ mod.Arithmetic.CN.I_in\[16\] _0638_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_50_216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5700_ _2116_ _2143_ _2145_ _2328_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_17_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6680_ mod.Data_Mem.F_M.dest\[8\] _3233_ _3234_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__3975__A2 mod.Arithmetic.CN.I_in\[32\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_1168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6889__I mod.Data_Mem.F_M.MRAM\[4\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5631_ _1840_ _2264_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5177__A1 _1745_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8350_ _0446_ net1 mod.Data_Mem.F_M.MRAM\[780\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5562_ _1542_ _2201_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__5972__I0 mod.Data_Mem.F_M.MRAM\[14\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7301_ _3617_ _0365_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4513_ _1090_ _1185_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_144_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_8281_ _0377_ net1 mod.Data_Mem.F_M.MRAM\[771\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5493_ _1690_ _2138_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_89_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7232_ _3576_ _0337_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__8234__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6221__S0 _2588_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6677__A1 mod.Data_Mem.F_M.dest\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4444_ _0928_ _1113_ _1115_ _1116_ _1117_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_99_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7163_ _3508_ mod.Data_Mem.F_M.MRAM\[12\]\[5\] _3534_ _3536_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4375_ _0968_ _0965_ _1048_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_98_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6429__A1 _2620_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6114_ mod.Data_Mem.F_M.MRAM\[1\]\[0\] _1539_ _1809_ mod.Data_Mem.F_M.MRAM\[0\]\[0\]
+ _2708_ _2731_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XTAP_430 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_59_817 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_7094_ mod.Data_Mem.F_M.MRAM\[23\]\[2\] _3494_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_100_402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_936 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8384__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6045_ mod.Data_Mem.F_M.MRAM\[16\]\[7\] mod.Data_Mem.F_M.MRAM\[17\]\[7\] _2540_ _2663_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_58_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5101__A1 _1764_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5033__I _1676_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3009 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7229__I0 _3523_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_820 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2308 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5968__I _1685_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2319 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_1046 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7996_ mod.P2.dest_reg1\[2\] net2 net1 mod.P2.dest_reg\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_42_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1607 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5404__A2 _1553_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1618 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1629 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6947_ _3405_ mod.Data_Mem.F_M.MRAM\[14\]\[7\] _3400_ _3406_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__4093__B _0748_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5955__A3 _2573_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_149_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_50_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6878_ _3361_ _0198_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_70_1208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5829_ mod.Data_Mem.F_M.MRAM\[18\]\[1\] mod.Data_Mem.F_M.MRAM\[19\]\[1\] _2452_ _2453_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_72_1090 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8548_ _0052_ net1 mod.Data_Mem.F_M.out_data\[28\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__6117__B1 _1575_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_159_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_163_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_8479_ _0575_ net1 mod.Data_Mem.F_M.MRAM\[797\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_135_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_1148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_151_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5652__B _2217_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4143__A2 _0818_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_430 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7468__I0 _3638_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5891__A2 mod.Data_Mem.F_M.MRAM\[771\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_134_52 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5878__I _2499_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2820 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2831 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2842 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2853 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5246__I2 _1907_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_503 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2864 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_17_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8107__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2875 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_127_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_32_216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2886 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2897 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_159_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_9_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5159__A1 _1804_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6356__B1 _2201_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8257__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_1204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7534__S _3745_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4134__A2 _0809_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5882__A2 _2501_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4160_ _0821_ _0835_ _0836_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_67_102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4091_ mod.Arithmetic.ACTI.x\[2\] _0768_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_23_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_820 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7850_ _3927_ _0603_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_75_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_503 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6801_ _3317_ _0165_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_36_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4993_ _1639_ _1661_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_7781_ _3887_ _0575_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_51_525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_95_1090 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6732_ _3234_ _3270_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__3948__A2 _0625_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3944_ _0621_ _0622_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6663_ mod.Data_Mem.F_M.MRAM\[27\]\[3\] _3222_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_104_1017 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5614_ mod.Data_Mem.F_M.MRAM\[797\]\[6\] _2226_ _1749_ mod.Data_Mem.F_M.MRAM\[796\]\[6\]
+ _2248_ _2249_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XANTENNA__6412__I _3020_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8402_ _0498_ net1 mod.Data_Mem.F_M.MRAM\[787\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_118_800 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6594_ _3187_ _0088_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_8333_ _0429_ net1 mod.Data_Mem.F_M.MRAM\[777\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__5570__A1 _2178_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5545_ _1533_ _2185_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_145_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_8264_ _0360_ net1 mod.Data_Mem.F_M.MRAM\[768\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5476_ _2074_ _2118_ _2119_ _2121_ _2123_ _0033_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_132_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7215_ _3531_ mod.Data_Mem.F_M.MRAM\[2\]\[3\] _3562_ _3566_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__4125__A2 _0670_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4427_ _1097_ _1098_ _1099_ _1100_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__4867__I _1535_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8195_ _0080_ net2 net1 mod.I_addr\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XANTENNA__6370__I0 _2032_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_1181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_120_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7146_ _3269_ _3270_ _3374_ _3524_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_4358_ _0627_ _1031_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4920__I1 mod.Data_Mem.F_M.MRAM\[768\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4088__B _0661_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_154_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_63_1056 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7077_ _3485_ _0273_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_47_809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_978 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4289_ _0960_ _0961_ _0957_ _0963_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_86_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6028_ _1670_ _2118_ _2639_ _2646_ _2647_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_39_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5698__I _1517_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2105 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_66_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2116 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2127 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_64_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_2138 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2149 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1404 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_588 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5389__A1 _1918_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_823 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1426 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_536 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7979_ _0205_ net1 mod.Data_Mem.F_M.MRAM\[4\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1437 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1448 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6050__A2 mod.Data_Mem.F_M.MRAM\[18\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1459 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_569 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_878 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_1152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4061__A1 _0674_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_168_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_74_1196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3946__I _0623_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4364__A2 _1024_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_135_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5313__A1 mod.Data_Mem.F_M.MRAM\[31\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5164__I1 mod.Data_Mem.F_M.MRAM\[786\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7153__I _3242_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6510__B1 _3110_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_145_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_133_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5616__A2 mod.Data_Mem.F_M.MRAM\[31\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5401__I _2061_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7613__I0 _3771_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2650 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2661 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2672 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2683 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2694 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1960 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_166_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1971 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1982 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1993 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6329__B1 _2157_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_158_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7328__I _3297_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5552__A1 mod.Data_Mem.F_M.MRAM\[29\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5330_ mod.Data_Mem.F_M.MRAM\[31\]\[6\] _1886_ _1993_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_154_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_114_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_115_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_1018 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5261_ mod.Data_Mem.F_M.MRAM\[799\]\[4\] _1913_ _1925_ _1926_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_48_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7000_ _3397_ mod.Data_Mem.F_M.MRAM\[17\]\[3\] _3435_ _3439_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4212_ _0825_ _0849_ _0887_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5192_ _1844_ _1857_ _1858_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_96_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4143_ _0802_ _0818_ _0819_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_96_753 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5607__A2 _2221_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_797 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4074_ mod.Arithmetic.CN.I_in\[17\] mod.Arithmetic.I_out\[73\] _0703_ _0751_ vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_83_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_680 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7902_ _0128_ net1 mod.Data_Mem.F_M.MRAM\[28\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_83_469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8422__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7833_ _0081_ _3917_ _0597_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_58_1136 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_169_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7764_ _3877_ _3878_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__4043__A1 _0710_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4976_ _1606_ _1644_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_11_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6715_ mod.Data_Mem.F_M.MRAM\[10\]\[0\] _3261_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__8572__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4594__A2 _1262_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7695_ _3841_ _0535_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5218__S1 _1882_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6646_ _3213_ _0114_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4346__A2 _0923_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6577_ mod.I_addr\[0\] mod.I_addr\[2\] mod.I_addr\[1\] _3176_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
X_8316_ _0412_ net1 mod.Data_Mem.F_M.MRAM\[775\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_133_611 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5528_ _1713_ _2169_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_30_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7296__A1 _1855_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8247_ _0343_ net1 mod.Data_Mem.F_M.MRAM\[30\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5459_ _2107_ _2108_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_105_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_160_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_132_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8178_ _0288_ net1 mod.Data_Mem.F_M.MRAM\[3\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_99_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7129_ _3514_ _0296_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_59_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_87_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_606 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_617 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_319 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_797 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4282__A1 _0806_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_1203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1201 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1212 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6559__B1 _3050_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6559__C2 _2496_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_163_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7349__S _3643_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1234 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_163_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_642 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_152_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_1245 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1256 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1267 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1278 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1289 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_539 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_109_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5385__I1 mod.Data_Mem.F_M.MRAM\[788\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_155_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_3_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_97_539 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7039__A1 _3464_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_1062 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5840__B _2463_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_904 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5332__S _1892_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8445__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_1213 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6262__A2 _1880_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3170 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3181 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3192 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8595__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7259__S _3590_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2480 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4830_ _1495_ _1499_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_2491 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_34_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4025__A1 mod.Arithmetic.CN.I_in\[23\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4761_ _1285_ _1323_ _1430_ _1431_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_53_1033 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1790 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1093 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_159_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6500_ _3083_ mod.Data_Mem.F_M.MRAM\[768\]\[4\] _3105_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_7480_ _3618_ mod.Data_Mem.F_M.MRAM\[780\]\[6\] _3713_ _3716_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_14_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4692_ _1350_ _1362_ _1363_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_6431_ _1536_ _3033_ _3035_ _3038_ _3039_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_6362_ _2868_ _2964_ _2972_ _2973_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_155_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5313_ mod.Data_Mem.F_M.MRAM\[31\]\[5\] _1759_ _1977_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_8101_ mod.Data_Mem.F_M.out_data\[11\] net2 net1 mod.Arithmetic.CN.I_in\[11\] vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_6293_ _2904_ mod.Data_Mem.F_M.MRAM\[15\]\[4\] mod.Data_Mem.F_M.MRAM\[14\]\[4\] _2905_
+ _2906_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_142_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6486__C1 _2502_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8032_ _0241_ net1 mod.Data_Mem.F_M.MRAM\[17\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5244_ mod.Data_Mem.F_M.MRAM\[771\]\[4\] mod.Data_Mem.F_M.MRAM\[770\]\[4\] _1908_
+ _1909_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_114_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_1184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5175_ _1835_ mod.Data_Mem.F_M.MRAM\[774\]\[3\] _1841_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__5242__S _1906_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4126_ _0631_ _0648_ _0802_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_84_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_907 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4057_ _0723_ _0728_ _0729_ _0733_ _0734_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_83_255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5976__I _2381_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7169__S _3534_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_642 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_169_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_36_193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4880__I _1504_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7816_ _3906_ _0591_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XPHY_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_51_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__7962__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_339 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_169_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6800__I1 _3316_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7747_ _3868_ _0560_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4959_ _1539_ _1627_ _1628_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_71_1144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_1155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7993__RN net2 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7678_ mod.Data_Mem.F_M.MRAM\[791\]\[7\] _3833_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_138_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_71_1199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8318__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6629_ mod.Data_Mem.F_M.MRAM\[26\]\[2\] _3205_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_137_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_106_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5216__I _1607_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8468__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_161_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_79_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_133_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8170__RN net2 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_904 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6492__A2 mod.Data_Mem.F_M.MRAM\[0\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_977 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_120_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_101_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_87_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_75_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4991__S _1658_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_90_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1020 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1042 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1053 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_16_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7744__A2 _3232_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1075 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_169_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1086 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5755__A1 _2187_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7984__RN net2 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5507__A1 _2138_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5327__S _1877_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_87_1162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7542__S _3752_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4030__I mod.Arithmetic.CN.I_in\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_83_1059 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4965__I _1616_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_859 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8161__RN net2 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7341__I _3635_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4494__A1 _1052_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5997__S _2331_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6235__A2 _1827_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_609 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6980_ _3397_ mod.Data_Mem.F_M.MRAM\[16\]\[3\] _3423_ _3427_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_81_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7985__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4097__I1 _0721_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5294__I0 mod.Data_Mem.F_M.MRAM\[771\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_65_288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5931_ _2548_ _2550_ _2551_ _2552_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_65_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5994__A1 _2587_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_1133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_642 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_146_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5862_ mod.Data_Mem.F_M.MRAM\[4\]\[2\] mod.Data_Mem.F_M.MRAM\[5\]\[2\] mod.Data_Mem.F_M.MRAM\[20\]\[2\]
+ mod.Data_Mem.F_M.MRAM\[21\]\[2\] _2025_ _2106_ _2485_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_33_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_1019 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7601_ _3765_ mod.Data_Mem.F_M.MRAM\[786\]\[3\] _3787_ _3792_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4813_ _1399_ _1474_ _1482_ _1483_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
X_8581_ _0597_ net1 mod.Instr_Mem.instruction\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5793_ _1675_ _2417_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_21_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7532_ _3748_ _0465_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4744_ _0622_ _1413_ _1414_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_30_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7463_ _3297_ _3705_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4675_ _1329_ _1345_ _1346_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_6414_ _2495_ _3023_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6171__A1 _1645_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_931 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7394_ _3670_ _0405_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6345_ _1608_ _1989_ _2763_ _2956_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__5036__I _1573_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_130_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6276_ _2846_ _2887_ _2888_ _2889_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_115_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8015_ _0224_ net1 mod.Data_Mem.F_M.MRAM\[15\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5227_ _1790_ _1892_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_88_358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6474__A2 _2304_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8152__RN net2 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_57_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5158_ _1805_ _1807_ _1810_ _1823_ _1824_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_29_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4109_ mod.Arithmetic.ACTI.x\[5\] _0786_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_72_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5089_ _1499_ _1756_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4237__A1 _0665_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4788__A2 _1344_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_72_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_114 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__5037__I0 _1702_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_125 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_136 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__8140__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_158 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_169_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_169 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_8_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4960__A2 _1628_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_166_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8290__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_739 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_10_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__8143__RN net2 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5899__S1 _1756_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6465__A2 _3069_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4476__A1 _1031_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_1081 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_121_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_169_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4228__A1 _0901_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_748 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_5 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_62_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5440__A3 _2076_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5028__I0 _1680_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_995 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4453__C mod.Arithmetic.ACTI.x\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_169_680 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7336__I _3305_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_156_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4460_ _1124_ _1132_ _1133_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__6153__A1 _2759_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4391_ _0843_ mod.Arithmetic.CN.I_in\[27\] _1064_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_139_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6130_ mod.Data_Mem.F_M.MRAM\[781\]\[1\] _2200_ _1809_ mod.Data_Mem.F_M.MRAM\[780\]\[1\]
+ _2746_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XTAP_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_645 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6061_ _2410_ _2674_ _2676_ _2678_ _2679_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XANTENNA__8134__RN net2 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8013__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_678 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5012_ _1675_ mod.Data_Mem.F_M.MRAM\[785\]\[1\] _1679_ _1680_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_66_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_1187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4219__A1 _0820_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_501 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6963_ _3252_ _3416_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__8163__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5914_ _2394_ _2535_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_146_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_50_910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6894_ _3369_ _0206_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_62_781 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_1015 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5845_ _2425_ mod.Data_Mem.F_M.MRAM\[785\]\[2\] _2468_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__3993__A3 _0669_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_166_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_10_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6351__S _2044_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8564_ _0068_ net1 mod.Data_Mem.F_M.out_data\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_33_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5776_ _2394_ _2099_ _2397_ _2400_ _2401_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_7515_ _3711_ mod.Data_Mem.F_M.MRAM\[782\]\[3\] _3734_ _3738_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_108_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4727_ _1282_ _1387_ _1397_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_8495_ _0591_ net1 mod.Data_Mem.F_M.MRAM\[7\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__4942__A2 _1610_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_148_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_717 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7446_ _3696_ _0431_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6144__A1 _2360_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6144__B2 _2188_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4658_ _1208_ _1207_ _1328_ _1217_ _1329_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_107_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7377_ mod.Data_Mem.F_M.MRAM\[773\]\[5\] _3662_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4589_ _1039_ _1144_ _1147_ _1261_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_103_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6328_ _2752_ _2939_ _2940_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_89_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8125__RN net2 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6447__A2 _2292_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6259_ _1663_ _2872_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_103_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_57_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8506__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6080__B1 mod.Data_Mem.F_M.MRAM\[15\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_718 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_461 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4630__A1 _1169_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_160_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_987 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6383__B2 _2992_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7156__I _3245_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_10_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_99_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_154_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_113_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8036__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4697__A1 _1134_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_84_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_68_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8116__RN net2 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4449__A1 _1007_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5110__A2 _1774_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8186__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7238__I1 mod.Data_Mem.F_M.MRAM\[30\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5340__S _1836_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_832 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5949__A1 _2567_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4464__B _1136_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3960_ _0636_ _0637_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4621__A1 _0731_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_1125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_1109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_148_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5630_ _2075_ _2263_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6374__A1 _2891_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4224__I1 _0897_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5561_ _1538_ _2200_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__5972__I1 mod.Data_Mem.F_M.MRAM\[15\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7300_ _3569_ mod.Data_Mem.F_M.MRAM\[768\]\[5\] _3608_ _3617_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4512_ _1169_ _1183_ _1184_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__6126__A1 _2366_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_536 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5492_ _2135_ mod.Data_Mem.F_M.MRAM\[30\]\[4\] _2136_ _2137_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_8280_ _0376_ net1 mod.Data_Mem.F_M.MRAM\[771\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_7231_ _3527_ mod.Data_Mem.F_M.MRAM\[30\]\[1\] _3574_ _3576_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__6221__S1 _2449_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_160_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4443_ _0915_ mod.Arithmetic.CN.I_in\[52\] _1116_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_99_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7162_ _3535_ _0308_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4374_ _0970_ _0974_ _1047_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_113_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_1216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8529__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6113_ _2728_ mod.Data_Mem.F_M.MRAM\[3\]\[0\] _1805_ _2729_ _2730_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XTAP_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8107__RN net2 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7093_ _3493_ _0281_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_101_915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_464 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6044_ _2379_ _2654_ _2661_ _2662_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__5101__A2 _1767_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_497 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_67_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7229__I1 mod.Data_Mem.F_M.MRAM\[30\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4860__A1 _1501_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2309 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7995_ mod.P2.dest_reg1\[1\] net2 net1 mod.P2.dest_reg\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_26_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1608 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6145__I _1573_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1619 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6946_ _3258_ _3405_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_169_17 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6877_ mod.Data_Mem.F_M.MRAM\[6\]\[6\] _3361_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_167_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5828_ _1519_ _2452_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__6365__A1 _2876_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8547_ _0051_ net1 mod.Data_Mem.F_M.out_data\[27\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_124_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5759_ mod.Data_Mem.F_M.MRAM\[782\]\[0\] mod.Data_Mem.F_M.MRAM\[783\]\[0\] _2383_
+ _2384_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_154_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_33_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8059__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_536 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8478_ _0574_ net1 mod.Data_Mem.F_M.MRAM\[797\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_108_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7429_ mod.Data_Mem.F_M.MRAM\[776\]\[7\] _3688_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_123_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6912__I0 _3249_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_150_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_89_464 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4446__A4 _1114_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_1212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_726 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_45_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_843 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2810 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2821 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2832 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2843 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2854 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2865 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2876 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2887 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_32_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2898 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_40_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6356__A1 mod.Data_Mem.F_M.MRAM\[13\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6356__B2 mod.Data_Mem.F_M.MRAM\[12\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_1180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6108__A1 _1640_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_1216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_153_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_355 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6903__I0 _3228_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_1082 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5619__B1 mod.Data_Mem.F_M.MRAM\[798\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4090_ _0749_ _0708_ _0762_ _0767_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_110_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4973__I _1529_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_501 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6800_ mod.Data_Mem.F_M.MRAM\[799\]\[5\] _3316_ _3313_ _3317_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_7780_ _3784_ mod.Data_Mem.F_M.MRAM\[797\]\[7\] _3883_ _3887_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4992_ _1608_ _1659_ _1614_ _1660_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_56_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6731_ _3231_ _3269_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_3943_ _0620_ _0621_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_56_1053 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4922__B _1590_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6662_ _3221_ _0122_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__8201__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6347__A1 _2012_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_31_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8401_ _0497_ net1 mod.Data_Mem.F_M.MRAM\[787\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_165_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5613_ _1940_ _2247_ _2248_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_136_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6593_ mod.Data_Mem.F_M.MRAM\[11\]\[0\] _3187_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_136_119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8332_ _0428_ net1 mod.Data_Mem.F_M.MRAM\[777\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_118_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_117_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5544_ _1804_ _2184_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_129_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5570__A2 _2199_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8351__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8263_ _0359_ net1 mod.Data_Mem.F_M.MRAM\[5\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5475_ _2095_ _2122_ _2123_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_117_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7214_ _3565_ _0330_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__7919__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4426_ _0833_ _1097_ _1099_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_8194_ net191 net2 net1 mod.Arithmetic.CN.F_in\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_8_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7145_ _3227_ _3523_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_67_1193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4357_ _0629_ _1028_ _1030_ mod.P3.Res\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_59_615 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_59_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7076_ mod.Data_Mem.F_M.MRAM\[21\]\[1\] _3485_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4288_ _0957_ _0960_ _0961_ _0962_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or3_1
XANTENNA__5086__A1 _1751_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_607 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_98_1109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4883__I _1551_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6027_ _2416_ _2641_ _2645_ _2646_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_104_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2106 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2117 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_640 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2128 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6035__B1 _2652_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2139 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1405 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1416 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4046__C1 _0721_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7978_ _0204_ net1 mod.Data_Mem.F_M.MRAM\[4\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1427 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1438 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1449 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6929_ _3393_ mod.Data_Mem.F_M.MRAM\[14\]\[1\] _3391_ _3394_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_126_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6338__A1 _1941_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_50_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5219__I _1653_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_155_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_6_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5849__B1 _2469_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_151_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__6510__A1 _1966_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5313__A2 _1759_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_924 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7310__I0 _3603_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5077__A1 _1742_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5889__I _1707_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_927 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_938 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_1020 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_161_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_18_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2640 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2651 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8224__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_1086 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2662 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_526 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2673 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2684 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5838__B _1804_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2695 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1950 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_159_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4052__A2 _0721_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1961 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1972 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1983 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6329__A1 mod.Data_Mem.F_M.MRAM\[781\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1994 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6329__B2 mod.Data_Mem.F_M.MRAM\[780\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_147_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8374__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4033__I _0709_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5552__A2 _1539_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4968__I _1594_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7829__A1 _3174_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_1084 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5260_ _1917_ _1924_ _1674_ _1925_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_141_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_114_358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_4211_ _0867_ _0885_ _0886_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_5191_ _1836_ mod.Data_Mem.F_M.MRAM\[769\]\[3\] _1856_ _1857_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_96_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_1208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4142_ _0812_ _0817_ _0818_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_95_220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5799__I _2422_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_765 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4073_ _0710_ _0750_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_49_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_95_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5863__I0 mod.Data_Mem.F_M.MRAM\[2\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7901_ _0127_ net1 mod.Data_Mem.F_M.MRAM\[27\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_3_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_83_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_48_191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7832_ _3916_ _3917_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_64_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_1148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7763_ _3230_ _3705_ _3371_ _3877_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_51_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4975_ mod.Data_Mem.F_M.MRAM\[6\]\[1\] _1640_ _1642_ _1643_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_6714_ _3260_ _0135_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6423__I _2388_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7694_ mod.Data_Mem.F_M.MRAM\[792\]\[7\] _3841_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6645_ mod.Data_Mem.F_M.MRAM\[25\]\[2\] _3213_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5039__I _1567_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_34_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6576_ _3174_ _3175_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__5543__A2 _2179_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4346__A3 _0840_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_164_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8315_ _0411_ net1 mod.Data_Mem.F_M.MRAM\[775\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_117_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5527_ _2132_ _2168_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_133_645 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8246_ _0342_ net1 mod.Data_Mem.F_M.MRAM\[30\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5458_ _2106_ _2107_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_117_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7891__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4409_ _1078_ _1081_ _1082_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_8177_ mod.P1.instr_reg\[8\] net2 net1 mod.P2.Rout_reg1\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_99_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5389_ _1918_ _2049_ _2050_ _2051_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_8_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7128_ _3445_ mod.Data_Mem.F_M.MRAM\[19\]\[0\] _3513_ _3514_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_115_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7059_ _3476_ _0264_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__8247__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4282__A2 mod.Arithmetic.CN.I_in\[19\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_1215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6559__A1 _3005_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1213 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6559__B2 _2652_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1224 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1235 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5658__B _2268_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8397__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1246 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1257 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3957__I _0633_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1268 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1279 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_30_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_168_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5534__A2 _2168_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5393__B _1775_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7531__I0 _3747_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_430 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5298__A1 _1633_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_112_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_1090 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5840__C _1498_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5412__I _2070_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_65_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_74_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_18_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3160 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_278 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3171 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_81 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3182 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3193 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2470 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5568__B _1631_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2481 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5222__A1 mod.Data_Mem.F_M.MRAM\[31\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2492 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6270__I0 _1895_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4760_ _1286_ _1322_ _1430_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_1780 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6970__A1 mod.Data_Mem.F_M.dest\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1791 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_53_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4691_ _1352_ _1361_ _1362_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_119_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_1078 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_1089 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6430_ _2560_ _2437_ _3037_ _2388_ _3038_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_146_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_127_461 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6361_ _2867_ _2971_ _2972_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_8100_ mod.Data_Mem.F_M.out_data\[10\] net2 net1 mod.Arithmetic.CN.I_in\[10\] vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_5312_ _1622_ _1975_ _1863_ _1976_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_6292_ _1493_ _2905_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__7522__I0 _3729_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6486__B1 _3030_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8031_ _0240_ net1 mod.Data_Mem.F_M.MRAM\[17\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_115_678 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5243_ _1587_ _1908_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__6486__C2 _2672_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_1163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5174_ _1690_ _1840_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_64_1196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4125_ _0649_ _0670_ _0801_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_84_713 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4056_ _0732_ _0733_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_83_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7815_ mod.Data_Mem.F_M.MRAM\[7\]\[7\] _3906_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XPHY_307 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_52_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_169_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__4016__A2 _0691_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_52_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7746_ _3771_ mod.Data_Mem.F_M.MRAM\[796\]\[0\] _3867_ _3868_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4958_ _1626_ _1627_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_123_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5992__I _2560_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7677_ _3832_ _0526_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_71_1167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4889_ _1557_ _1558_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6628_ _3204_ _0105_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4319__A3 _0838_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7761__I0 _3784_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_165_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6559_ _3005_ _2350_ _3050_ _2652_ _2650_ _2496_ _3161_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_106_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7513__I0 _3640_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_106_678 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_160_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_121_615 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8229_ mod.P1.instr_reg\[11\] net2 net1 mod.P2.dest_reg1\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_0_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_121_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_31 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5827__I0 mod.Data_Mem.F_M.MRAM\[2\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_746 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1010 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1021 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1032 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_35_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5204__A1 _1802_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1054 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_71_985 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7744__A3 _3634_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1065 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_71_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1087 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_169_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_7_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6180__A2 _2200_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4191__A1 _0812_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8412__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_152_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_1174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_805 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7622__I _3801_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_816 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_83_1049 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_151_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5691__A1 _2319_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4494__A2 _1074_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8562__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5294__I1 mod.Data_Mem.F_M.MRAM\[770\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5930_ _2512_ mod.Data_Mem.F_M.MRAM\[773\]\[4\] _2551_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_59_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5861_ _2416_ _2473_ _2483_ _2484_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_34_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_90_1009 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7600_ _1787_ _3789_ _3791_ _0490_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_61_473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4812_ _1477_ _1479_ _1481_ _1482_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_21_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8580_ _0596_ net1 mod.Instr_Mem.instruction\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__5746__A2 _2364_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5792_ _2378_ _2416_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_159_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7531_ _3747_ mod.Data_Mem.F_M.MRAM\[783\]\[1\] _3745_ _3748_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4743_ mod.Arithmetic.CN.I_in\[47\] _1412_ _1413_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__4954__B1 _1621_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7462_ _3704_ _0439_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_119_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4674_ _1234_ _1344_ _1345_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_147_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6413_ mod.Data_Mem.F_M.MRAM\[0\]\[0\] mod.Data_Mem.F_M.MRAM\[1\]\[0\] _2258_ _3022_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__5903__C1 _2524_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7393_ mod.Data_Mem.F_M.MRAM\[774\]\[5\] _3670_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6171__A2 _1680_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8092__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6344_ _1635_ _1990_ _2955_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_1_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_131_913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_153_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6275_ _2872_ _1905_ _2888_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_103_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8014_ _0223_ net1 mod.Data_Mem.F_M.MRAM\[14\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5226_ mod.Data_Mem.F_M.MRAM\[21\]\[4\] mod.Data_Mem.F_M.MRAM\[20\]\[4\] _1890_ _1891_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_131_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_69_540 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4377__B _0877_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4485__A2 _1141_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5157_ _1653_ _1815_ _1821_ _1822_ _1823_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_57_746 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4108_ _0735_ _0778_ _0784_ _0785_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_5088_ _1508_ _1741_ _1754_ _1755_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_38_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_57_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5434__A1 _2080_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_278 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_112_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_429 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4039_ _0715_ _0716_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_71_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_749 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7187__A1 _3294_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_974 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_80_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__5037__I1 _1703_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_126 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_148 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_169_158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_36_1040 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_7729_ _3858_ _0552_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_40_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5936__B _2100_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_1084 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_138_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__8435__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_1213 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5227__I _1790_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4131__I _0806_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_106_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8585__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_161_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_133_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5673__A1 _2288_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_797 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_75_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_532 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5425__A1 _2081_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3987__A1 _0633_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_6 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_16_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5028__I1 _1684_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_646 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_1140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4936__B1 _1603_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7617__I _3797_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__4400__A2 _1072_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_157_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_12_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4041__I mod.Arithmetic.I_out\[72\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4164__A1 _0617_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4390_ _1062_ _1063_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_98_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__8595__D _0611_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4976__I _1606_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7952__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6060_ _2565_ _2677_ _2678_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__6456__A3 _3062_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_646 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4467__A2 _1122_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5011_ _1677_ _1678_ _1679_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_39_724 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_1155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_852 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8308__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_1199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4219__A2 _0826_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_513 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6962_ _3415_ _0228_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_53_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5913_ _1726_ _2534_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_6893_ mod.Data_Mem.F_M.MRAM\[4\]\[6\] _3369_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_22_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_62_771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4216__I _0653_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8458__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_793 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5844_ _2464_ _2466_ _2467_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_34_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8563_ _0067_ net1 mod.Data_Mem.F_M.out_data\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5775_ _2313_ mod.Data_Mem.F_M.MRAM\[788\]\[0\] _2399_ _2400_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__6392__A2 _2993_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7514_ _3737_ _0458_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4726_ _1276_ _1388_ _1389_ _1273_ _1396_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_120_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_8494_ _0590_ net1 mod.Data_Mem.F_M.MRAM\[7\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_7445_ mod.Data_Mem.F_M.MRAM\[777\]\[7\] _3696_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6144__A2 mod.Data_Mem.F_M.MRAM\[6\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4657_ _1206_ _1212_ _1328_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5047__I _1646_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4155__A1 _0655_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7376_ _3661_ _0396_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4588_ _1149_ _1152_ _1259_ _1260_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_104_913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_162_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6327_ _2904_ mod.Data_Mem.F_M.MRAM\[783\]\[5\] mod.Data_Mem.F_M.MRAM\[782\]\[5\]
+ _2267_ _2939_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_143_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_88_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6258_ _2870_ _1874_ _2871_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_66_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5655__A1 _2091_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5209_ mod.Data_Mem.F_M.MRAM\[5\]\[4\] mod.Data_Mem.F_M.MRAM\[4\]\[4\] _1873_ _1874_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_6189_ _2360_ mod.Data_Mem.F_M.MRAM\[6\]\[2\] mod.Data_Mem.F_M.MRAM\[7\]\[2\] _2188_
+ _2804_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_29_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_690 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_532 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5510__I _1779_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_546 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6080__A1 _2696_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3969__A1 _0645_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6080__B2 _2517_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4630__A2 _1183_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_41_977 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4570__B _0634_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3965__I _0641_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_166_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4997__S _1636_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4146__A1 _0652_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7975__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_1111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5894__A1 _2511_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_84_1155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_1188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4449__A2 _1015_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_513 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5420__I _1489_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5949__A2 mod.Data_Mem.F_M.MRAM\[2\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_63_546 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6071__A1 _2172_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_169_1087 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4036__I _0702_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_793 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_1148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6374__A2 _2040_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5068__S _1658_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4385__A1 _0616_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5560_ mod.Data_Mem.F_M.MRAM\[797\]\[2\] _2179_ _2195_ mod.Data_Mem.F_M.MRAM\[796\]\[2\]
+ _2198_ _2199_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XFILLER_129_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_117_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4511_ _1058_ _1172_ _1182_ _1183_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_156_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_526 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5491_ _1791_ mod.Data_Mem.F_M.MRAM\[31\]\[4\] _2136_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__6126__A2 _2195_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_1055 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7230_ _3575_ _0336_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4442_ mod.Arithmetic.CN.I_in\[50\] _1114_ _1115_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_89_1088 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5885__A1 _2266_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7161_ _3533_ mod.Data_Mem.F_M.MRAM\[12\]\[4\] _3534_ _3535_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4373_ _1044_ _1045_ _1046_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_98_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6112_ _2540_ mod.Data_Mem.F_M.MRAM\[2\]\[0\] _2729_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XTAP_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_7092_ mod.Data_Mem.F_M.MRAM\[23\]\[1\] _3493_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_432 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8130__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_465 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6043_ _2434_ _2660_ _2661_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_498 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4860__A2 _1528_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7994_ mod.P2.dest_reg1\[0\] net2 net1 mod.P2.dest_reg\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XANTENNA__8280__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6062__A1 _2531_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1609 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6945_ _3404_ _0222_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_81_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4612__A2 _1187_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_730 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6876_ _3360_ _0197_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_5827_ mod.Data_Mem.F_M.MRAM\[2\]\[1\] mod.Data_Mem.F_M.MRAM\[3\]\[1\] _1954_ _2451_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_10_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_50_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6365__A2 _2024_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_796 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4376__A1 _0966_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7998__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5758_ _1588_ _2383_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_8546_ _0050_ net1 mod.Data_Mem.F_M.out_data\[26\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_148_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4709_ _1373_ _1379_ _1380_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__6117__A2 _1505_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8477_ _0573_ net1 mod.Data_Mem.F_M.MRAM\[797\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__7314__A1 _3610_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5689_ _2312_ _2137_ _2314_ _2317_ _2318_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_159_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7428_ _3687_ _0422_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6912__I1 mod.Data_Mem.F_M.MRAM\[13\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5876__A1 _2496_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7359_ mod.Data_Mem.F_M.MRAM\[772\]\[4\] _3653_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_78_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_103_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_131_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5628__A1 _2089_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_32 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_131_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_100_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2800 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_17_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_57_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2811 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_166_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_150_31 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2822 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6053__A1 _2185_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2833 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2844 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2855 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2866 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4603__A2 _1258_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2877 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2888 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2899 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_129_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_752 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_40_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_1110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__8003__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_159_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_90_1192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_167_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_154_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6903__I1 mod.Data_Mem.F_M.MRAM\[13\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8153__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_890 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6020__B _2638_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_1061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5415__I _2073_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_49_1094 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_68_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_150_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_48_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6044__A1 _2379_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4991_ mod.Data_Mem.F_M.MRAM\[19\]\[1\] mod.Data_Mem.F_M.MRAM\[18\]\[1\] _1658_ _1659_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__4055__B1 _0730_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6730_ _3268_ _0143_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_56_1021 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_398 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3942_ _0619_ _0620_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_32_730 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_output7_I net7 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_6661_ mod.Data_Mem.F_M.MRAM\[27\]\[2\] _3221_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6347__A2 _1988_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5612_ _2233_ mod.Data_Mem.F_M.MRAM\[799\]\[6\] mod.Data_Mem.F_M.MRAM\[798\]\[6\]
+ _2234_ _2247_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
X_8400_ _0496_ net1 mod.Data_Mem.F_M.MRAM\[787\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_158_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6592_ _3186_ _0087_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_30_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_8331_ _0427_ net1 mod.Data_Mem.F_M.MRAM\[777\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5543_ mod.Data_Mem.F_M.MRAM\[797\]\[1\] _2179_ _1640_ mod.Data_Mem.F_M.MRAM\[796\]\[1\]
+ _2182_ _2183_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XFILLER_157_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8262_ _0358_ net1 mod.Data_Mem.F_M.MRAM\[5\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5474_ mod.Data_Mem.F_M.MRAM\[798\]\[1\] mod.Data_Mem.F_M.MRAM\[799\]\[1\] _1908_
+ _2122_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_160_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5858__A1 _2440_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7213_ _3529_ mod.Data_Mem.F_M.MRAM\[2\]\[2\] _3562_ _3565_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4425_ _0619_ mod.Arithmetic.CN.I_in\[41\] _0897_ _0984_ _1098_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_8193_ _0303_ net1 mod.Data_Mem.F_M.MRAM\[19\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_99_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7144_ _3522_ _0303_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4356_ _0775_ _0855_ _0856_ _1029_ _0627_ _1030_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_98_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_584 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7075_ _3484_ _0272_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_59_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_284 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4287_ _0915_ _0959_ _0808_ _0873_ _0961_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XFILLER_86_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_969 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_100_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6026_ _2642_ _2643_ _2644_ _2565_ _2645_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_101_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2107 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6035__A1 _2539_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2118 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2129 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6035__B2 _2435_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1406 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7977_ _0203_ net1 mod.Data_Mem.F_M.MRAM\[4\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_42_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1417 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1428 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1439 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8026__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4597__A1 mod.Arithmetic.ACTI.x\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6928_ _3239_ _3393_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_167_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_161_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6859_ mod.Data_Mem.F_M.MRAM\[779\]\[5\] _3352_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_35_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_11_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6338__A2 _2002_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4349__A1 _0992_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8176__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_149_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8529_ _0033_ net1 mod.Data_Mem.F_M.out_data\[41\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__5149__I0 mod.Data_Mem.F_M.MRAM\[3\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_159_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5849__B2 _2403_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_104_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_893 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_104_584 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6267__S _2723_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_1169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5171__S _1836_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5077__A2 _1743_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6274__A1 _1941_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_822 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_1032 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6026__A1 _2642_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6026__B2 _2565_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2630 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_166_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2641 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6577__A2 mod.I_addr\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2652 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2663 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2674 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_398 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4588__A1 _1149_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2685 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1940 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1951 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2696 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1962 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1973 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8519__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1984 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6329__A2 _2751_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1995 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_103_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_1052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_155_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_103_1096 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__7561__S _3760_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5145__I _1503_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4210_ _0881_ _0884_ _0885_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__4512__A1 _1169_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5190_ _1658_ _1855_ _1856_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_69_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4141_ _0815_ _0816_ _0817_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_96_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4072_ _0675_ _0705_ _0749_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_55_107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6360__S1 _2750_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7900_ _0126_ net1 mod.Data_Mem.F_M.MRAM\[27\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__5863__I1 mod.Data_Mem.F_M.MRAM\[3\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8049__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6905__S _3376_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xtiny_user_project_170 wbs_dat_o[23] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XANTENNA__6017__A1 _2061_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7831_ _0612_ _3175_ _3916_ _0596_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_91_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_1029 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6704__I _3252_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4974_ _1641_ _1642_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_7762_ _3876_ _0567_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_51_335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5776__B1 _2397_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8199__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6713_ _3259_ mod.Data_Mem.F_M.MRAM\[28\]\[7\] _3250_ _3260_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_149_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7693_ _3840_ _0534_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_165_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6644_ _3212_ _0113_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5379__I0 mod.Data_Mem.F_M.MRAM\[771\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8517__185 net185 vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
X_6575_ mod.I_addr\[3\] _3174_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_30_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_1212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8314_ _0410_ net1 mod.Data_Mem.F_M.MRAM\[775\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5526_ _2081_ _2067_ _2159_ _2165_ _2166_ _2167_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XANTENNA__4751__A1 _1203_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_118_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_161_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8245_ _0341_ net1 mod.Data_Mem.F_M.MRAM\[30\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_133_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5457_ _1495_ _2106_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_105_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4408_ _0716_ _0816_ _0972_ _1080_ _1081_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
X_8176_ mod.P1.instr_reg\[7\] net2 net1 mod.P2.Rout_reg1\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_5388_ _1875_ mod.Data_Mem.F_M.MRAM\[786\]\[7\] _2050_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_120_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7127_ _3512_ _3513_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_113_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4894__I _1562_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4339_ _1010_ _1012_ _1013_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_87_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_532 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7058_ mod.Data_Mem.F_M.MRAM\[20\]\[0\] _3476_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_47_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_1191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6009_ _2104_ _2627_ _2628_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_27_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_55_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7056__I0 _3462_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1203 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6559__A2 _2350_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1214 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1225 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1236 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1247 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1258 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1269 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5862__S0 _2025_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_128_429 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_168_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_155_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3973__I _0645_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5534__A3 _2174_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5166__S _1581_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4070__S _0746_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4742__A1 _1411_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_151_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6495__A1 _2353_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7531__I1 mod.Data_Mem.F_M.MRAM\[783\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_722 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7039__A3 _3335_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_497 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6247__A1 _2107_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_1045 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_38_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_78_788 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3150 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3161 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_34_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3172 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8341__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_994 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3183 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8228__RN net2 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3194 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2460 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2471 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7909__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2482 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2493 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5222__A2 _1886_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6270__I1 _1893_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1770 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1062 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1781 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1792 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_147_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8491__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_390 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4690_ _1359_ _1360_ _1361_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__4979__I _1646_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7355__I mod.Data_Mem.F_M.MRAM\[772\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5076__S _1519_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4733__A1 mod.Arithmetic.CN.I_in\[61\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6360_ _2246_ _2249_ _2967_ _2970_ _1964_ _2750_ _2971_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_143_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5311_ _1969_ _1970_ _1973_ _1974_ _1695_ _1795_ _1975_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_114_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6291_ _2059_ _2904_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__7522__I1 mod.Data_Mem.F_M.MRAM\[782\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8030_ _0239_ net1 mod.Data_Mem.F_M.MRAM\[16\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__6486__A1 _3026_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5242_ mod.Data_Mem.F_M.MRAM\[769\]\[4\] mod.Data_Mem.F_M.MRAM\[768\]\[4\] _1906_
+ _1907_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__6486__B2 _2497_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5173_ _1828_ _1831_ _1833_ _1838_ _1839_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__7090__I mod.Data_Mem.F_M.MRAM\[23\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6238__A1 _2160_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4124_ _0629_ _0671_ _0800_ mod.P3.Res\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_60_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_69_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xinput1 io_in[8] net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_20
XFILLER_84_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4055_ _0725_ _0727_ _0730_ _0731_ _0732_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_84_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_65_950 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_983 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7814_ _3905_ _0590_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_24_335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_290 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_319 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__6410__A1 _3017_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_169_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7745_ _3866_ _3867_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_4957_ _1501_ _1553_ _1626_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_51_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7466__S _3707_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6370__S _1738_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7676_ mod.Data_Mem.F_M.MRAM\[791\]\[6\] _3832_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4888_ _1556_ _1557_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_137_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_20_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_1179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4889__I _1557_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6627_ mod.Data_Mem.F_M.MRAM\[26\]\[1\] _3204_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_20_596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5367__I3 _2028_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7761__I1 mod.Data_Mem.F_M.MRAM\[796\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4724__A1 _0789_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6558_ _2353_ _2347_ _2663_ _2642_ _3159_ _3160_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_119_985 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5509_ _2144_ _2151_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_69_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_646 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6489_ _3082_ _3094_ _0075_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__8214__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8228_ mod.P1.instr_reg\[10\] net2 net1 mod.P2.dest_reg1\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_121_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_830 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_8159_ mod.Data_Mem.F_M.out_data\[69\] net2 net1 mod.Arithmetic.CN.I_in\[69\] vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XANTENNA__6229__A1 _2838_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8364__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4129__I _0804_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5988__B1 _2397_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5452__A2 _1554_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3968__I _0641_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1000 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_942 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1022 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_1046 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1033 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5204__A2 _1803_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6401__A1 _2418_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1055 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1066 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1077 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_169_852 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1088 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_129_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_169_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7201__I0 _3508_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7175__I mod.Data_Mem.F_M.MRAM\[22\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_52_1090 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_167_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_125_911 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_109_473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6468__A1 _3017_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_1077 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_1088 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_806 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_83_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_817 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_98_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_32_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_78_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_39_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5691__A2 mod.Data_Mem.F_M.MRAM\[797\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_427 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4039__I _0715_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_1200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_674 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6254__I _2702_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5860_ _2474_ _2482_ _2483_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_34_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_1108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_1157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_1119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5826__S0 _2025_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4811_ _1363_ _1383_ _1480_ _1481_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_2290 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_107_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_34_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5791_ _2415_ _0056_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__7881__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_61_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4742_ _1411_ mod.Arithmetic.CN.I_in\[46\] _1412_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_7530_ _3302_ _3747_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4954__A1 _1620_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4954__B2 mod.Data_Mem.F_M.MRAM\[783\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_7461_ mod.Data_Mem.F_M.MRAM\[778\]\[7\] _3704_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4673_ _1334_ _1343_ _1344_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__8237__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6412_ _3020_ _3021_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5903__B1 _2523_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7392_ _3669_ _0404_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_162_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6343_ _2882_ _2952_ _2953_ _2884_ _1898_ _2954_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_127_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_1204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6459__A1 _2619_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6274_ _1941_ _1904_ _2887_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_88_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8387__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8013_ _0222_ net1 mod.Data_Mem.F_M.MRAM\[14\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5225_ _1587_ _1890_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__5131__A1 _1759_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7259__I0 mod.Data_Mem.F_M.MRAM\[31\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5156_ _1530_ _1822_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_29_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_213 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4890__B1 mod.Data_Mem.F_M.MRAM\[31\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4107_ _0730_ _0778_ _0784_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5087_ _1744_ _1748_ _1750_ _1753_ _1616_ _1754_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_56_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5434__A2 _2077_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4038_ mod.Arithmetic.CN.I_in\[10\] _0715_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_84_588 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_430 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_964 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_169_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7187__A2 _3464_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_116 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_52_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5198__A1 mod.Data_Mem.F_M.MRAM\[783\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_127 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_25_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_5989_ _1620_ _2601_ _2602_ _2104_ _2378_ _2608_ _2609_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai222_1
XPHY_149 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6490__S0 _2290_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7728_ mod.Data_Mem.F_M.MRAM\[795\]\[0\] _3858_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5936__C _2449_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_166_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6113__B _1805_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7659_ _3823_ _0517_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_165_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_118_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_977 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_498 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5122__A1 _1714_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_1050 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_1061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5673__A2 mod.Data_Mem.F_M.MRAM\[28\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_1056 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_87_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_43_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_48_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5425__A2 _0010_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_739 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6074__I _2685_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_430 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3987__A2 mod.Arithmetic.ACTI.x\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_44_975 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6386__B1 _2201_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6802__I net9 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4936__A1 mod.Data_Mem.F_M.MRAM\[790\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_156_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_30_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_129_546 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5418__I _2076_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5736__I0 mod.Data_Mem.F_M.MRAM\[16\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5361__A1 mod.Data_Mem.F_M.MRAM\[15\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4164__A2 mod.Arithmetic.CN.I_in\[57\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7489__I0 _3638_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_936 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_603 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5113__A1 _1779_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_647 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5010_ mod.Data_Mem.F_M.MRAM\[784\]\[1\] _1678_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_1123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_500 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_39_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_1167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_38_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_717 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6961_ _3399_ _1870_ _3414_ _3415_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_93_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_1030 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_249 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5912_ _2080_ _2520_ _2533_ _0059_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_6892_ _3368_ _0205_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_59_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5843_ _2417_ _1787_ _2465_ _2466_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_61_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6712__I _3258_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4927__A1 _1595_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8562_ _0066_ net1 mod.Data_Mem.F_M.out_data\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_148_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_146_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5774_ _2398_ mod.Data_Mem.F_M.MRAM\[789\]\[0\] _2399_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_7513_ _3640_ mod.Data_Mem.F_M.MRAM\[782\]\[2\] _3734_ _3737_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4725_ _1272_ _1390_ _1395_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_8493_ _0589_ net1 mod.Data_Mem.F_M.MRAM\[7\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_147_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7444_ _3695_ _0430_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4656_ _1219_ _1325_ _1326_ _1327_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_163_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_730 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5352__A1 _1933_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4155__A2 mod.Arithmetic.CN.I_in\[41\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7375_ mod.Data_Mem.F_M.MRAM\[773\]\[4\] _3661_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_66_1001 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4587_ _1154_ _1158_ _1258_ _1259_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_118_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6326_ mod.Data_Mem.F_M.MRAM\[13\]\[5\] _2901_ _2902_ mod.Data_Mem.F_M.MRAM\[12\]\[5\]
+ _2937_ _2938_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XANTENNA__6159__I _2713_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5104__A1 _1708_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6257_ _1574_ _2870_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_77_809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_103_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5208_ _1587_ _1873_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__5655__A2 _1803_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6188_ _2798_ _2802_ _2703_ _2803_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_130_287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_680 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_393 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5139_ _1641_ _1805_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_57_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_897 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_739 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_1130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6080__A2 mod.Data_Mem.F_M.MRAM\[14\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_290 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3969__A2 mod.Arithmetic.CN.I_in\[24\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_569 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_1163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8402__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_603 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_1185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4570__C _0775_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_31 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_12_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__8552__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_126_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4146__A2 _0657_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_153_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_49_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5894__A2 _1846_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4697__A3 _1366_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_284 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6069__I _2685_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_1167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_755 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5902__S _2321_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6843__A1 _3316_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_801 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_739 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6018__B _2354_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6071__A2 _2687_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8082__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_249 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_867 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_355 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_761 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_143_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_157_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_31_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4385__A2 _0691_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5582__A1 _2211_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4510_ _1180_ _1181_ _1182_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_89_1023 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_1094 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5490_ _2134_ _2135_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_8_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_145_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4441_ _0616_ mod.Arithmetic.CN.I_in\[51\] _1114_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_7160_ _3524_ _3534_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_4372_ _0976_ _1024_ _1045_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6111_ _1691_ _2728_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_98_433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7091_ _3492_ _0280_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_59_809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_433 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_99_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6042_ _2423_ _2655_ _2656_ _2464_ _2659_ _2660_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_101_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6707__I net9 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8425__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_82_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_897 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_739 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7993_ mod.Instr_Mem.instruction\[30\] net2 net1 mod.Data_Mem.F_M.src\[8\] vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_6944_ _3403_ mod.Data_Mem.F_M.MRAM\[14\]\[6\] _3400_ _3404_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_82_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_81_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8575__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6875_ mod.Data_Mem.F_M.MRAM\[6\]\[5\] _3360_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_50_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6442__I _2499_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5826_ mod.Data_Mem.F_M.MRAM\[4\]\[1\] mod.Data_Mem.F_M.MRAM\[5\]\[1\] mod.Data_Mem.F_M.MRAM\[20\]\[1\]
+ mod.Data_Mem.F_M.MRAM\[21\]\[1\] _2025_ _2106_ _2450_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_23_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_22_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4376__A2 _0965_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8545_ _0049_ net1 mod.Data_Mem.F_M.out_data\[25\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5757_ _2381_ _2382_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5058__I _1725_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4708_ _1374_ _1378_ _1379_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_159_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8476_ _0572_ net1 mod.Data_Mem.F_M.MRAM\[797\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_108_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5688_ _2315_ mod.Data_Mem.F_M.MRAM\[28\]\[4\] _2316_ _2317_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__7314__A2 _3626_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4897__I _1565_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7427_ mod.Data_Mem.F_M.MRAM\[776\]\[6\] _3687_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_118_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4639_ _0844_ mod.Arithmetic.CN.I_in\[22\] _0678_ _1310_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_135_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5876__A2 _2497_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_162_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7358_ _3652_ _0387_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_89_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6309_ _1978_ _1979_ _2723_ _2921_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_104_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7289_ _3302_ _3610_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5628__A2 _2099_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_820 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_92_609 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5521__I _1812_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2801 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2812 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2823 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6053__A2 _2154_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2834 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4137__I _0637_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_168_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2845 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2856 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2867 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_32_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2878 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2889 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3976__I _0616_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7942__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4367__A2 _0974_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_13_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_166_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4119__A2 _0673_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_49_1051 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6020__C _2263_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8448__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5619__A2 mod.Data_Mem.F_M.MRAM\[799\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_714 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_71 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5431__I _1549_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_82_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7559__S _3760_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4047__I mod.Arithmetic.CN.I_in\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_64_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4990_ _1646_ _1658_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_23_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4055__B2 _0731_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_1000 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3941_ _0618_ _0619_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_56_1033 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_1055 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6660_ _3220_ _0121_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_5611_ mod.Data_Mem.F_M.MRAM\[29\]\[6\] _2086_ _2227_ mod.Data_Mem.F_M.MRAM\[28\]\[6\]
+ _2245_ _2246_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XFILLER_83_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5555__A1 _2178_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6591_ mod.I_addr\[7\] _3185_ _3186_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_129_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_8330_ _0426_ net1 mod.Data_Mem.F_M.MRAM\[777\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5542_ _2180_ _2181_ _2182_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_8_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_858 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8261_ _0357_ net1 mod.Data_Mem.F_M.MRAM\[5\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5473_ _2097_ mod.Data_Mem.F_M.MRAM\[30\]\[1\] _2120_ _2121_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_117_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7212_ _3564_ _0329_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4424_ _0897_ _0984_ _1097_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_144_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8192_ _0302_ net1 mod.Data_Mem.F_M.MRAM\[19\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_28_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_67_1162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_160_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_390 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7143_ _3462_ mod.Data_Mem.F_M.MRAM\[19\]\[7\] _3518_ _3522_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4355_ _0775_ _0774_ _0794_ _1029_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_63_1015 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7821__I _3910_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_63_1048 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7074_ mod.Data_Mem.F_M.MRAM\[21\]\[0\] _3484_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_58_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4286_ _0959_ _0808_ _0873_ _0960_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_100_202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_101_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6025_ mod.Data_Mem.F_M.MRAM\[14\]\[6\] mod.Data_Mem.F_M.MRAM\[15\]\[6\] _2360_ _2644_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_55_801 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7607__I0 _3782_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_95_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_536 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_171 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2108 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6035__A2 _2650_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2119 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_867 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7976_ _0202_ net1 mod.Data_Mem.F_M.MRAM\[4\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1407 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7965__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1418 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1429 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6927_ _3392_ _0216_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_42_539 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_74_1144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6858_ _3351_ _0188_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_168_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_74_1188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4349__A2 _1002_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5809_ _2421_ _2432_ _2433_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_6789_ net6 _3308_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_167_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_148_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8528_ _0032_ net1 mod.Data_Mem.F_M.out_data\[40\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_108_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5149__I1 mod.Data_Mem.F_M.MRAM\[1\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8459_ _0555_ net1 mod.Data_Mem.F_M.MRAM\[795\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__5516__I _1543_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5849__A2 _2125_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_163_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_1213 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_49_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6274__A2 _1904_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6026__A2 _2643_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_1055 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2620 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2631 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2642 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_675 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2653 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2664 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2675 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1930 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2686 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1941 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2697 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1952 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1963 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1974 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1985 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7526__A2 _3705_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1996 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_9_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8120__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6810__I mod.Data_Mem.F_M.MRAM\[789\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_167_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_1004 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4760__A2 _1322_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__8270__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_1048 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5870__B _1804_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4512__A2 _1183_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5362__S _1879_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4140_ _0621_ mod.Arithmetic.CN.I_in\[8\] _0709_ _0816_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XANTENNA__6257__I _1574_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4071_ mod.Arithmetic.ACTI.x\[1\] _0748_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_56_609 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_789 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7988__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_981 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_1100 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_1111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xtiny_user_project_160 wbs_dat_o[13] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_48_171 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtiny_user_project_171 wbs_dat_o[24] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_48_193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6017__A2 mod.Data_Mem.F_M.MRAM\[18\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_149_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7830_ _3915_ _3916_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4028__A1 _0674_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5076__I0 mod.Data_Mem.F_M.MRAM\[17\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7761_ _3784_ mod.Data_Mem.F_M.MRAM\[796\]\[7\] _3872_ _3876_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__5776__A1 _2394_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4973_ _1529_ _1641_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_52_859 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5776__B2 _2400_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6712_ _3258_ _3259_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_32_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7692_ mod.Data_Mem.F_M.MRAM\[792\]\[6\] _3840_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6643_ mod.Data_Mem.F_M.MRAM\[25\]\[1\] _3212_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5379__I1 mod.Data_Mem.F_M.MRAM\[770\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_149_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6574_ _3173_ _0082_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4200__A1 _0844_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_146_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8313_ _0409_ net1 mod.Data_Mem.F_M.MRAM\[775\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5525_ _2114_ _2166_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__4751__A2 mod.Arithmetic.CN.I_in\[46\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7752__S _3867_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4240__I _0807_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_156_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_117_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_8244_ _0340_ net1 mod.Data_Mem.F_M.MRAM\[30\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5456_ _2081_ _2104_ _2105_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_145_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4407_ _0715_ _0972_ _1079_ _1080_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_161_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8175_ mod.DM_en net2 net1 mod.DMen_reg vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XANTENNA__5700__A1 _2116_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5387_ mod.Data_Mem.F_M.MRAM\[787\]\[7\] _2049_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_132_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7126_ _3433_ _3407_ _3421_ _3512_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_59_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4338_ _0914_ _1011_ _1012_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_75_907 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7057_ _3475_ _0263_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_47_609 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4269_ _0862_ _0943_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__5071__I _1737_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6008_ mod.Data_Mem.F_M.MRAM\[770\]\[6\] mod.Data_Mem.F_M.MRAM\[771\]\[6\] _2275_
+ _2627_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__7199__S _3553_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7056__I1 mod.Data_Mem.F_M.MRAM\[1\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_15_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1204 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1215 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8143__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1226 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5767__A1 _2210_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_163_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7959_ _0185_ net1 mod.Data_Mem.F_M.MRAM\[779\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5311__S0 _1695_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1248 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1259 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5862__S1 _2106_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7996__RN net2 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_11_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_7_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8293__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_149_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6192__A1 _1742_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4742__A2 mod.Arithmetic.CN.I_in\[46\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_109_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8173__RN net2 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6495__A2 _3095_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_1081 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_46_1054 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_77_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_46_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4258__A1 _0929_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_20_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_93_759 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3140 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3151 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3162 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5849__C _2471_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3173 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3184 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3195 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2450 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2461 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2472 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2483 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2494 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6741__S _3274_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_1161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7987__RN net2 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1760 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1771 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1782 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_1025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1793 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6183__A1 _2206_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5230__I0 mod.Data_Mem.F_M.MRAM\[17\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5930__A1 _2512_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5156__I _1530_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4733__A2 _1366_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_161_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7572__S _3773_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4060__I mod.Arithmetic.CN.I_in\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_155_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5310_ mod.Data_Mem.F_M.MRAM\[3\]\[5\] mod.Data_Mem.F_M.MRAM\[2\]\[5\] _1968_ _1974_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_6290_ _1564_ _2903_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_127_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4995__I _1525_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6486__A2 _2309_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5241_ _1835_ _1906_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__8164__RN net2 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7371__I mod.Data_Mem.F_M.MRAM\[773\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8016__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5172_ _1834_ _1837_ _1838_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_96_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4123_ _0661_ _0796_ _0798_ _0799_ _0628_ _0800_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XANTENNA__6916__S _3381_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4249__A1 _0619_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_68_277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4054_ mod.Arithmetic.CN.I_in\[13\] _0731_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput2 io_in[9] net2 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_20
XFILLER_49_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8166__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7813_ mod.Data_Mem.F_M.MRAM\[7\]\[6\] _3905_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_64_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__6410__A2 mod.Data_Mem.F_M.MRAM\[13\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_7744_ _3230_ _3232_ _3634_ _3866_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_52_678 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4956_ _1489_ _1625_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_80_998 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7675_ _3831_ _0525_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_20_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4887_ _1553_ _1555_ _1556_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6626_ _3203_ _0104_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6174__A1 _1898_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5921__A1 _2097_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6557_ _2312_ _2508_ _2668_ _1757_ _3159_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_118_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_923 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_5508_ _2119_ _2148_ _2150_ _2133_ _0038_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
X_6488_ _3003_ _3091_ _3093_ _3094_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_156_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8227_ mod.P1.instr_reg\[9\] net2 net1 mod.P2.dest_reg1\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XANTENNA__8155__RN net2 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5439_ _2090_ _0025_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__7281__I _3292_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8158_ mod.Data_Mem.F_M.out_data\[68\] net2 net1 mod.Arithmetic.CN.I_in\[68\] vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_114_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_59_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8509__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7109_ _3502_ _0288_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_87_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_8089_ mod.P2.Rout_reg1\[1\] net2 net1 mod.P2.Rout_reg\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_102_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5988__A1 _2394_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5988__B2 _2604_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_718 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4660__A1 _0651_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_167_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1001 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1023 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1058 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_150_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1045 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1056 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_678 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4412__A1 _1002_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_169_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1078 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1089 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3984__I mod.Arithmetic.ACTI.x\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7201__I1 mod.Data_Mem.F_M.MRAM\[29\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_168_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6165__A1 _1706_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5912__A1 _2080_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8039__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5905__S _2331_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_124_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_1154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6468__A2 mod.Data_Mem.F_M.MRAM\[1\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8146__RN net2 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_1198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_680 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8189__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_4_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5979__A1 _2301_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4100__B1 _0774_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_962 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4651__A1 _1297_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_1125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7567__S _3759_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_1169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5826__S1 _2106_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2280 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_22_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4810_ _1365_ _1382_ _1480_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XTAP_2291 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_464 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5790_ _1491_ _2372_ _2374_ _2412_ _2414_ _2415_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai32_1
XANTENNA__4403__A1 _0893_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5600__B1 _1749_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1590 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4741_ _1338_ _1411_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_7460_ _3703_ _0438_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4672_ _1337_ _1341_ _1342_ _1343_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_31_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_1180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6411_ _2376_ _3020_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5903__A1 _2517_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4706__A2 _1376_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_761 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7391_ mod.Data_Mem.F_M.MRAM\[774\]\[4\] _3669_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6342_ _2015_ _2016_ _1738_ _2953_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_66_1216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6459__A2 mod.Data_Mem.F_M.MRAM\[0\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8137__RN net2 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6273_ _2686_ _2886_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_88_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8012_ _0221_ net1 mod.Data_Mem.F_M.MRAM\[14\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_102_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5224_ mod.Data_Mem.F_M.MRAM\[23\]\[4\] mod.Data_Mem.F_M.MRAM\[22\]\[4\] _1588_ _1889_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_29_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5131__A2 _1796_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7259__I1 _3316_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5155_ _1557_ _1818_ _1820_ _1821_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_69_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_575 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_726 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4890__A1 mod.Data_Mem.F_M.MRAM\[15\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4890__B2 _1558_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4106_ _0771_ _0777_ _0780_ _0781_ _0782_ _0783_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
X_5086_ _1751_ _1752_ _1753_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_84_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_759 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4037_ _0687_ _0683_ _0713_ _0714_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_84_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4642__A1 _1063_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7187__A3 _3335_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_106 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__6381__S _1881_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_117 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_128 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__5198__A2 _1863_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5988_ _2394_ _2142_ _2397_ _2604_ _2607_ _2608_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XPHY_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_52_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7727_ _3857_ _0551_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6490__S1 _2171_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4939_ _1607_ _1608_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_21_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7658_ mod.Data_Mem.F_M.MRAM\[790\]\[5\] _3823_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_20_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6609_ mod.Data_Mem.F_M.MRAM\[24\]\[0\] _3195_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_166_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_7589_ _3321_ _3784_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_119_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_21_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5952__C _2572_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_107_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_77 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8331__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8128__RN net2 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5122__A2 mod.Data_Mem.F_M.MRAM\[787\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_1035 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_501 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_788 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4881__A1 _1548_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8481__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_47_225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_759 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3979__I mod.Arithmetic.CN.I_in\[40\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_8 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_15_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_43_464 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_987 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6386__A1 mod.Data_Mem.F_M.MRAM\[13\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6386__B2 mod.Data_Mem.F_M.MRAM\[12\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_1120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4936__A2 _1601_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6304__B _2873_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_169_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_8_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_1164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6090__I _2706_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_1017 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6138__A1 _2752_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5736__I1 mod.Data_Mem.F_M.MRAM\[17\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5361__A2 _1886_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8119__RN net2 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_98_615 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_604 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_615 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_1113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5370__S _1588_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4872__A1 mod.Data_Mem.F_M.src\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7110__I0 _3450_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_1179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_320 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_504 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6960_ _3408_ _3414_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_5911_ _2526_ _2532_ _2533_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_4_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6891_ mod.Data_Mem.F_M.MRAM\[4\]\[5\] _3368_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_50_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8204__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6377__A1 _2872_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5842_ _2418_ mod.Data_Mem.F_M.MRAM\[787\]\[2\] _2465_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_107_1007 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_1220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8561_ _0065_ net1 mod.Data_Mem.F_M.out_data\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5773_ _1658_ _2398_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_22_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_166_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4513__I _1090_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7512_ _3736_ _0457_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4724_ _0789_ _1266_ _1268_ _1394_ mod.P3.Res\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__6129__A1 _2619_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8492_ _0588_ net1 mod.Data_Mem.F_M.MRAM\[7\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__6129__B2 _2089_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7443_ mod.Data_Mem.F_M.MRAM\[777\]\[6\] _3695_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__8354__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_148_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4655_ _1222_ _1256_ _1326_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_107_219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_162_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_539 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7374_ _3660_ _0395_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5352__A2 _2013_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4586_ _1197_ _1201_ _1257_ _1258_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XANTENNA__7629__A1 _2013_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_1013 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6325_ _2903_ _2936_ _2937_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_104_915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_1057 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6256_ _2686_ _2869_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5104__A2 _1770_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5207_ _1550_ _1872_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6187_ _2687_ _2801_ _1965_ _2802_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_5138_ _1799_ _1804_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_85_843 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5069_ _1734_ _1735_ _1736_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_44_217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4615__A1 _1205_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6108__C _2715_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_773 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7000__S _3435_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_1197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_968 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5519__I _1527_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_165_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_154_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6540__A1 _2619_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_797 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7871__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6843__A2 _3337_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_501 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4854__A1 _1522_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_88_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_48_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_169_1001 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_36_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_48_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_95 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8227__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_773 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6359__A1 mod.Data_Mem.F_M.MRAM\[781\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6359__B2 mod.Data_Mem.F_M.MRAM\[780\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8377__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_148_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5429__I _1725_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4385__A3 mod.Arithmetic.CN.I_in\[19\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5582__A2 _2212_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_1051 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7859__A1 _3913_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_5 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5365__S _1877_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4440_ mod.Arithmetic.CN.I_in\[52\] _0997_ _1113_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__6531__A1 _3106_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_160_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_132_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_99_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4371_ _0978_ _1043_ _1044_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_113_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6110_ _2185_ _2717_ _2726_ _2727_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XTAP_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7090_ mod.Data_Mem.F_M.MRAM\[23\]\[0\] _3492_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7331__I0 _3603_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_434 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6041_ _2548_ _2657_ _2658_ _2659_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XTAP_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_86_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_467 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6390__S0 _1489_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_67_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7992_ mod.Instr_Mem.instruction\[26\] net2 net1 mod.Data_Mem.F_M.src\[4\] vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_93_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_96_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6943_ _3255_ _3403_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_54_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6062__A3 _2679_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6874_ _3359_ _0196_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_50_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5825_ _2448_ _2449_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_167_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_72_1050 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8544_ _0048_ net1 mod.Data_Mem.F_M.out_data\[24\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5756_ _2380_ _2381_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_147_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_4707_ _1375_ _1377_ _1378_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_136_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_8475_ _0571_ net1 mod.Data_Mem.F_M.MRAM\[797\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5687_ _2267_ _2316_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_108_539 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_163_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7426_ _3686_ _0421_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6522__A1 _2321_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4638_ _1180_ _1308_ _1309_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__7894__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7357_ mod.Data_Mem.F_M.MRAM\[772\]\[3\] _3652_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4569_ _0614_ mod.Arithmetic.CN.I_in\[69\] _1241_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_104_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6308_ _2869_ _2919_ _2920_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_103_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7322__I0 _3569_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7288_ _3608_ _3609_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6286__B1 _2897_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_789 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6239_ _2846_ _2851_ _2852_ _2853_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__4836__A1 _1501_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_40_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_962 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6834__S _3337_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2802 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2813 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2824 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2835 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2846 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2857 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4064__A2 _0740_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5261__A1 mod.Data_Mem.F_M.MRAM\[799\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2868 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2879 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_159_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5249__I _1503_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_1161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5693__B _2311_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_86_1208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7561__I0 _3725_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6513__A1 _2528_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_153_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_142_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_4_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5712__I _2025_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5875__I0 mod.Data_Mem.F_M.MRAM\[786\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_759 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_898 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_751 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4055__A2 _0727_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5252__A1 _1700_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_51_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3940_ _0617_ _0618_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_90_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_149_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5610_ _2228_ _2244_ _2245_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_31_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6590_ _3178_ mod.I_addr\[6\] mod.I_addr\[5\] _3179_ _3185_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XANTENNA__5555__A2 _2183_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5541_ _1782_ mod.Data_Mem.F_M.MRAM\[799\]\[1\] mod.Data_Mem.F_M.MRAM\[798\]\[1\]
+ _2009_ _2181_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_118_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5095__S _1746_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_145_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8260_ _0356_ net1 mod.Data_Mem.F_M.MRAM\[5\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5472_ _1951_ mod.Data_Mem.F_M.MRAM\[31\]\[1\] _2120_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_7211_ _3527_ mod.Data_Mem.F_M.MRAM\[2\]\[1\] _3562_ _3564_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4423_ _0654_ mod.Arithmetic.CN.I_in\[44\] _1096_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_8191_ _0301_ net1 mod.Data_Mem.F_M.MRAM\[19\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_132_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_7142_ _3521_ _0302_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4354_ _0942_ _1027_ _1028_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_63_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_1185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_607 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7073_ _3483_ _0271_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4285_ _0958_ _0959_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_87_949 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4818__A1 _0673_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6024_ mod.Data_Mem.F_M.MRAM\[2\]\[6\] mod.Data_Mem.F_M.MRAM\[3\]\[6\] _2528_ _2643_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_86_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_651 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_95_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8542__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5491__A1 _1791_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4294__A2 _0966_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7607__I1 mod.Data_Mem.F_M.MRAM\[786\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2109 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7975_ _0201_ net1 mod.Data_Mem.F_M.MRAM\[4\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_81_131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4046__A2 _0708_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1408 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6453__I _2499_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6440__B1 _3046_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6926_ _3386_ mod.Data_Mem.F_M.MRAM\[14\]\[0\] _3391_ _3392_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_35_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6857_ mod.Data_Mem.F_M.MRAM\[779\]\[4\] _3351_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_74_1167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5808_ _2423_ _2122_ _2427_ _2403_ _2431_ _2432_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_22_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4349__A3 _1022_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6788_ _3307_ _0162_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_109_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8527_ net179 net1 mod.Data_Mem.F_M.out_data\[55\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5739_ mod.Data_Mem.F_M.MRAM\[4\]\[0\] mod.Data_Mem.F_M.MRAM\[5\]\[0\] mod.Data_Mem.F_M.MRAM\[20\]\[0\]
+ mod.Data_Mem.F_M.MRAM\[21\]\[0\] _1714_ _1756_ _2364_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__7284__I _3605_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8458_ _0554_ net1 mod.Data_Mem.F_M.MRAM\[795\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__5149__I2 mod.Data_Mem.F_M.MRAM\[0\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7409_ mod.Data_Mem.F_M.MRAM\[775\]\[5\] _3678_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_8389_ _0485_ net1 mod.Data_Mem.F_M.MRAM\[785\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_123_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8072__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_145_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4809__A1 _1372_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5482__A1 _2110_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4148__I _0620_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_610 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2610 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2621 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2632 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5234__A1 _1898_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2643 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2654 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2665 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1920 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2676 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1931 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1942 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2687 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2698 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1953 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1964 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1975 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1986 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1997 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_158_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_9_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_16_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8415__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7534__I0 _3749_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6498__B1 _2536_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6739__S _3274_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_391 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4767__B _1422_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8565__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_96_724 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_110_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4070_ _0630_ _0704_ _0746_ _0747_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__5473__A1 _2097_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4058__I _0731_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xtiny_user_project_150 wbs_dat_o[3] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_161 wbs_dat_o[14] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_3_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_49_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_1123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xtiny_user_project_172 wbs_dat_o[25] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_63_120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7369__I mod.Data_Mem.F_M.MRAM\[773\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_1129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6273__I _2686_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7760_ _3875_ _0566_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_36_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4972_ _1639_ _1640_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_17_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5776__A2 _2099_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6711_ net10 _3258_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5110__C _1508_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7691_ _3839_ _0533_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6025__I0 mod.Data_Mem.F_M.MRAM\[14\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6642_ _3211_ _0112_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_32_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6573_ _3171_ _3172_ _3173_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_160_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__4200__A2 mod.Arithmetic.CN.I_in\[18\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8140__D mod.Data_Mem.F_M.out_data\[50\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8095__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8312_ _0408_ net1 mod.Data_Mem.F_M.MRAM\[775\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_69_1203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5524_ mod.Data_Mem.F_M.MRAM\[29\]\[0\] _2087_ _2160_ _2164_ _2165_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_118_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4751__A3 _1208_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_106_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_8243_ _0339_ net1 mod.Data_Mem.F_M.MRAM\[30\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5455_ _2100_ _2103_ _2104_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__7832__I _3916_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4406_ _0813_ _0722_ _0715_ mod.Arithmetic.CN.I_in\[9\] _1079_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
X_8174_ mod.P2.dest_reg\[8\] net2 net1 mod.Data_Mem.F_M.dest\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_160_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5386_ _1700_ _2047_ _2048_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5700__A2 _2143_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7125_ _3511_ _0295_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_59_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4337_ _0641_ mod.Arithmetic.ACTI.x\[3\] _1011_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_99_584 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7932__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7056_ _3462_ mod.Data_Mem.F_M.MRAM\[1\]\[7\] _3465_ _3475_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4268_ _0861_ _0938_ _0942_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_68_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6007_ _1757_ _2626_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_74_429 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4199_ mod.Arithmetic.CN.I_in\[24\] _0809_ _0873_ _0874_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_67_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_1207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7279__I mod.Data_Mem.F_M.MRAM\[5\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_816 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_83_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1216 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7958_ _0184_ net1 mod.Data_Mem.F_M.MRAM\[779\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1227 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5311__S1 _1795_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5767__A2 _2387_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1238 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_646 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1249 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6909_ _3246_ mod.Data_Mem.F_M.MRAM\[13\]\[3\] _3376_ _3380_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_70_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7889_ _0115_ net1 mod.Data_Mem.F_M.MRAM\[25\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_168_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6911__I _3375_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8438__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_13_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6192__A2 _1739_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_164_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__8588__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5463__S _1873_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_163_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_152_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_104_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5262__I _1653_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_1014 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_1066 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5455__A1 _2100_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_77_278 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3130 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3141 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3152 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3163 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_3174 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6404__B1 _2384_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2440 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3185 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_3196 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2451 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2462 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2473 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2484 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2495 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1750 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4966__B1 _1633_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1761 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1772 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1783 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1794 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7755__I0 _3778_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_159_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5437__I _2088_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6183__A2 _2682_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5230__I1 mod.Data_Mem.F_M.MRAM\[16\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4194__A1 _0644_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_154_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5373__S _1894_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7955__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5240_ mod.Data_Mem.F_M.MRAM\[775\]\[4\] mod.Data_Mem.F_M.MRAM\[774\]\[4\] _1836_
+ _1905_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_142_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5694__A1 _2280_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5171_ mod.Data_Mem.F_M.MRAM\[789\]\[3\] mod.Data_Mem.F_M.MRAM\[788\]\[3\] _1836_
+ _1837_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_116_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_1155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_746 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_843 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4122_ _0794_ _0799_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_96_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_57_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_1188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5446__A1 _2091_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4249__A2 mod.Arithmetic.CN.I_in\[57\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_429 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4053_ _0679_ _0698_ _0713_ _0730_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_83_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5900__I _1609_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6932__S _3391_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7812_ _3904_ _0589_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_52_646 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7743_ _3865_ _0559_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_80_988 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4955_ _1618_ _1623_ _1624_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_162_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4421__A2 _1093_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7674_ mod.Data_Mem.F_M.MRAM\[791\]\[5\] _3831_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_60_690 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7746__I0 _3771_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4886_ _1554_ _1537_ _1555_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_32_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_1159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6625_ mod.Data_Mem.F_M.MRAM\[26\]\[0\] _3203_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6174__A2 _2789_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_146_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6556_ _3021_ _2677_ _3157_ _2108_ _3158_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XANTENNA__5921__A2 mod.Data_Mem.F_M.MRAM\[786\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5507_ _2138_ mod.Data_Mem.F_M.MRAM\[798\]\[6\] _2149_ _2150_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_3_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6487_ _3004_ _3092_ _3093_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_145_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8226_ _0327_ net1 mod.Data_Mem.F_M.MRAM\[29\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5438_ _2089_ _2067_ _2090_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_82_1200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_161_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5685__A1 _2313_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8157_ mod.Data_Mem.F_M.out_data\[67\] net2 net1 mod.Arithmetic.CN.I_in\[67\] vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XANTENNA__5082__I _1600_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5369_ mod.Data_Mem.F_M.MRAM\[31\]\[7\] _1913_ _2031_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_43_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_832 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7108_ _3445_ mod.Data_Mem.F_M.MRAM\[3\]\[0\] _3501_ _3502_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_59_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8088_ mod.P2.Rout_reg1\[0\] net2 net1 mod.P2.Rout_reg\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_87_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8110__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_23 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_87_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7039_ _3464_ _3332_ _3335_ _3465_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_59_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5988__A2 _2142_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5810__I _2100_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7003__S _3440_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3999__A1 _0674_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_462 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_985 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_911 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4660__A2 mod.Arithmetic.CN.I_in\[35\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1002 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1013 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8260__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6398__C1 _2404_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1035 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1046 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1057 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1068 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4412__A2 _1022_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8091__RN net2 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_24_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_7_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7978__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5912__A2 _2520_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_124_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7472__I _3308_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_819 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_151_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_105_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_34_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4651__A2 _1300_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_47_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6752__S _3279_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_61_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_1137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_146_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_34_646 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6779__I1 _3293_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2270 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2281 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2292 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_21_307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5600__A1 mod.Data_Mem.F_M.MRAM\[797\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4403__A2 _0829_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5600__B2 mod.Data_Mem.F_M.MRAM\[796\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4740_ _1407_ _1409_ _1410_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_1591 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4671_ _1338_ _1209_ _1342_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_30_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6410_ _3017_ mod.Data_Mem.F_M.MRAM\[13\]\[0\] _2382_ _3018_ _3019_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__4071__I mod.Arithmetic.ACTI.x\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7390_ _3668_ _0403_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5903__A2 _2521_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_1192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6341_ mod.Data_Mem.F_M.MRAM\[789\]\[6\] mod.Data_Mem.F_M.MRAM\[791\]\[6\] mod.Data_Mem.F_M.MRAM\[790\]\[6\]
+ mod.Data_Mem.F_M.MRAM\[788\]\[6\] _2448_ _1932_ _2952_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_155_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_127_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6272_ _2880_ _2882_ _2883_ _2884_ _1490_ _2885_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_143_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_153_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_130_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8011_ _0220_ net1 mod.Data_Mem.F_M.MRAM\[14\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__8133__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5223_ _1550_ _1888_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_69_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_532 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_69_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5154_ _1584_ _1819_ _1820_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_57_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5419__A1 _2072_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4105_ _0776_ _0774_ _0782_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__4890__A2 _1536_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5085_ mod.Data_Mem.F_M.MRAM\[21\]\[2\] mod.Data_Mem.F_M.MRAM\[20\]\[2\] _1701_ _1752_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_110_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5630__I _2075_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8283__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6092__A1 _1764_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_1048 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_1059 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4036_ _0702_ _0713_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_72_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_911 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_53_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_793 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_966 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_107 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__5786__B _2410_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5987_ _2406_ _2605_ _2606_ _2403_ _2607_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XPHY_118 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8073__RN net2 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_129 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_169_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_796 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7726_ mod.Data_Mem.F_M.MRAM\[794\]\[7\] _3857_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4938_ _1606_ _1607_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_75_1081 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4869_ _1537_ _1538_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_7657_ _3822_ _0516_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_162_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7493__S _3720_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6608_ _3194_ _0095_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_7588_ _3783_ _0486_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_20_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_118_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6539_ _2522_ mod.Data_Mem.F_M.MRAM\[781\]\[6\] _3142_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__6410__B _2382_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7292__I _3305_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5805__I _2395_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5658__A1 _2288_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8209_ _0310_ net1 mod.Data_Mem.F_M.MRAM\[12\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_133_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6837__S _3340_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_1052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4330__A1 _0921_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_82_1085 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_153_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4881__A2 _1549_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_169_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6083__A1 _1802_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_31 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_43_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_9 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_43_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3995__I mod.P2.Rout_reg\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6386__A2 _1538_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_785 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_796 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8006__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_1132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_85 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_169_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_168_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_11_362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4149__A1 _0824_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5897__A1 _2416_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8156__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_156_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_109_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_426 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4321__A1 _0654_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_1125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4872__A2 _1503_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_568 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7578__S _3773_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5821__A1 _2434_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_1021 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5910_ _2457_ _2530_ _2531_ _1800_ _2532_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_46_270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6890_ _3367_ _0204_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_62_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5841_ _2109_ _2464_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_146_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_785 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_1019 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_498 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5772_ _2396_ _2397_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_8560_ _0064_ net1 mod.Data_Mem.F_M.out_data\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_21_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4723_ _1031_ _1392_ _1393_ _1394_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_7511_ _3638_ mod.Data_Mem.F_M.MRAM\[782\]\[1\] _3734_ _3736_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_8491_ _0587_ net1 mod.Data_Mem.F_M.MRAM\[7\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__6129__A2 mod.Data_Mem.F_M.MRAM\[783\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7442_ _3694_ _0429_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4654_ _1222_ _1256_ _1325_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_107_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7373_ mod.Data_Mem.F_M.MRAM\[773\]\[3\] _3660_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4935__I0 mod.Data_Mem.F_M.MRAM\[789\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4585_ _1219_ _1222_ _1256_ _1257_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XANTENNA__5625__I _1845_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6324_ _2134_ mod.Data_Mem.F_M.MRAM\[15\]\[5\] mod.Data_Mem.F_M.MRAM\[14\]\[5\] _2905_
+ _2936_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_157_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6688__I0 _3240_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_724 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_104_949 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6255_ _2867_ _2868_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_89_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6301__A2 _2900_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5206_ _1870_ _1673_ _1871_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_88_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_800 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6186_ mod.Data_Mem.F_M.MRAM\[13\]\[2\] _2200_ _2202_ mod.Data_Mem.F_M.MRAM\[12\]\[2\]
+ _2800_ _2801_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_130_278 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5137_ _1669_ _1626_ _1803_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5360__I _2022_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5068_ mod.Data_Mem.F_M.MRAM\[1\]\[2\] mod.Data_Mem.F_M.MRAM\[0\]\[2\] _1658_ _1735_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_45_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_57_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5812__A1 _2152_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8029__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4019_ _0695_ _0696_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_16_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_53_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7287__I _3605_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4379__A1 _0687_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8179__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_7709_ _3848_ _0542_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_21_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5736__S _2360_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_166_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_138_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6540__A2 mod.Data_Mem.F_M.MRAM\[780\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_49_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4551__A1 _0929_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_84_1125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_162_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4303__A1 _0927_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_800 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6056__A1 _2672_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_169_1013 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4067__B1 _0740_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_1180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5803__A1 _2424_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_169_1068 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_90_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6359__A2 _2751_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_785 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7556__A1 _3612_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5567__B1 _2202_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_498 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_169_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5582__A3 _2219_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7859__A2 _3917_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6531__A2 mod.Data_Mem.F_M.MRAM\[13\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4542__A1 _0636_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4370_ _0990_ _1023_ _1043_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_99_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_936 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_63_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_402 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_152_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5381__S _1908_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6295__A1 mod.Data_Mem.F_M.MRAM\[13\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6295__B2 mod.Data_Mem.F_M.MRAM\[12\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6040_ _2549_ mod.Data_Mem.F_M.MRAM\[772\]\[7\] _2658_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_86_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_65_1080 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_800 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_67_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_468 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6390__S1 _2750_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_121_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_66_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6047__A1 _2214_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_27_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_1007 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7991_ mod.Instr_Mem.instruction\[24\] net2 net1 mod.Data_Mem.F_M.src\[2\] vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_54_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_1018 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_538 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6942_ _3402_ _0221_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_81_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8321__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6873_ mod.Data_Mem.F_M.MRAM\[6\]\[4\] _3359_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_23_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_22_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5824_ _2234_ _2448_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_50_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8543_ _0047_ net1 mod.Data_Mem.F_M.out_data\[39\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5755_ _2187_ _2064_ _2380_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_120_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__8471__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4706_ _1241_ _1376_ _1377_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_108_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6507__C1 _2541_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5686_ _1675_ _2315_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_8474_ _0570_ net1 mod.Data_Mem.F_M.MRAM\[797\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_148_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_162_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7425_ mod.Data_Mem.F_M.MRAM\[776\]\[5\] _3686_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4637_ _0633_ _0958_ _1062_ _1307_ _1308_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_68_1109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8200__RN net2 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6522__A2 mod.Data_Mem.F_M.MRAM\[768\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7771__S _3878_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4533__A1 _1203_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7356_ _3651_ _0386_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4533__B2 _1095_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4568_ _1238_ _1131_ _1239_ _1240_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_2_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_150_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_29 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6307_ _2915_ _2916_ _2917_ _2918_ _2919_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_7287_ _3605_ _3608_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__7322__I1 mod.Data_Mem.F_M.MRAM\[770\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4499_ _1055_ _1064_ _1070_ _1171_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_103_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5333__I0 mod.Data_Mem.F_M.MRAM\[19\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6238_ _2160_ _1842_ _2852_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_83_1191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4836__A2 _1504_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5090__I _1756_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_980 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6169_ _2186_ _1694_ _2785_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_1216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2803 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_23 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2814 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2825 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2836 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2847 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2858 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2869 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_25_251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6210__A1 _2196_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7745__I _3866_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_1184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_167_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_126_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6513__A2 mod.Data_Mem.F_M.MRAM\[0\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5265__I _1929_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7561__I1 mod.Data_Mem.F_M.MRAM\[784\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_1091 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_134_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_49_1086 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6277__A1 _1826_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5324__I0 mod.Data_Mem.F_M.MRAM\[5\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_939 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4827__A2 _1495_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5875__I1 mod.Data_Mem.F_M.MRAM\[787\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8344__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_611 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5252__A2 _1916_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_677 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_891 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4344__I _1017_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_1046 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8494__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_290 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__4763__A1 _1251_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5540_ _1572_ _2180_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_144_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5471_ _2090_ _2119_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_69_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_7210_ _3563_ _0328_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4422_ _1091_ _1094_ _1095_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_160_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_8190_ _0300_ net1 mod.Data_Mem.F_M.MRAM\[19\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_126_871 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7141_ _3460_ mod.Data_Mem.F_M.MRAM\[19\]\[6\] _3518_ _3521_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_119_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4353_ _0945_ _1026_ _1027_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_99_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_1197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7072_ mod.Data_Mem.F_M.MRAM\[20\]\[7\] _3483_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_59_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4284_ mod.Arithmetic.CN.I_in\[27\] _0958_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_86_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4818__A2 _0674_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_427 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6023_ _2388_ _2642_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6935__S _3391_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_67_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5491__A2 mod.Data_Mem.F_M.MRAM\[31\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7974_ _0200_ net1 mod.Data_Mem.F_M.MRAM\[4\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_81_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1409 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6440__A1 _3030_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6440__B2 _2672_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6925_ _3390_ _3391_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_74_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_63_891 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6856_ _3350_ _0187_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_22_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7240__I0 _3569_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_167_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_161_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5807_ _2428_ _1687_ _2429_ _2430_ _2431_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_3999_ _0674_ mod.Arithmetic.I_out\[79\] _0675_ _0676_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XANTENNA__5286__S _1612_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6787_ mod.Data_Mem.F_M.MRAM\[799\]\[2\] _3306_ _3300_ _3307_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_22_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4754__A1 _1185_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8526_ net180 net1 mod.Data_Mem.F_M.out_data\[54\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5738_ _2112_ _2355_ _2357_ _2359_ _2361_ _2362_ _2363_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_136_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_149_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_163_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8457_ _0553_ net1 mod.Data_Mem.F_M.MRAM\[795\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5669_ _2074_ _2118_ _2293_ _2299_ _0050_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_135_134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8217__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7408_ _3677_ _0412_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_159_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_8388_ _0484_ net1 mod.Data_Mem.F_M.MRAM\[785\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_85_1220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_151_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7339_ _3531_ mod.Data_Mem.F_M.MRAM\[771\]\[3\] _3636_ _3642_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_116_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_939 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8367__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_104_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4809__A2 _1380_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6845__S _3340_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5482__A2 _2127_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_1013 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_161_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_782 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2600 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2611 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2622 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2633 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5234__A2 _1628_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6431__A1 _1536_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2644 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_31 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1910 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2655 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2666 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1921 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2677 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1932 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2688 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_72_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1943 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_159_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2699 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1954 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1965 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1976 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7231__I0 _3527_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1987 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1998 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4745__A1 _0622_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_155_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_85 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_126_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7534__I1 mod.Data_Mem.F_M.MRAM\[783\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6498__A1 _2353_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_1088 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6498__B2 _2556_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_114_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_830 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4767__C mod.Arithmetic.ACTI.x\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7298__I0 _3615_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_69_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_427 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_1050 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5473__A2 mod.Data_Mem.F_M.MRAM\[30\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_1083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xtiny_user_project_140 la_data_out[61] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_64_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
Xtiny_user_project_151 wbs_dat_o[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_23_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xtiny_user_project_162 wbs_dat_o[15] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_37_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xtiny_user_project_173 wbs_dat_o[26] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_92_942 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7470__I0 _3640_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4971_ _1600_ _1639_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__7884__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6710_ _3257_ _0134_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4984__A1 _1645_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7690_ mod.Data_Mem.F_M.MRAM\[792\]\[5\] _3839_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA_output5_I net5 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6025__I1 mod.Data_Mem.F_M.MRAM\[15\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_149_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6641_ mod.Data_Mem.F_M.MRAM\[25\]\[0\] _3211_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6186__B1 _2202_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6503__B _3107_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_73_1190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4736__A1 _1293_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6572_ _0612_ _3169_ _3172_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_8311_ _0407_ net1 mod.Data_Mem.F_M.MRAM\[774\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_145_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5523_ _2163_ _2164_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__5834__S _2398_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8242_ _0338_ net1 mod.Data_Mem.F_M.MRAM\[30\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5454_ _2102_ _2103_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_161_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_133_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_132_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_4405_ _0620_ _0724_ _1078_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_8173_ mod.P2.dest_reg\[4\] net2 net1 mod.Data_Mem.F_M.dest\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_5385_ mod.Data_Mem.F_M.MRAM\[791\]\[7\] mod.Data_Mem.F_M.MRAM\[788\]\[7\] mod.Data_Mem.F_M.MRAM\[789\]\[7\]
+ mod.Data_Mem.F_M.MRAM\[790\]\[7\] _1829_ _2009_ _2047_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__5633__I _1875_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5700__A3 _2145_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_1051 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7124_ _3462_ mod.Data_Mem.F_M.MRAM\[3\]\[7\] _3506_ _3511_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4336_ _0642_ mod.Arithmetic.ACTI.x\[2\] _0842_ _1010_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_59_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7055_ _3474_ _0262_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_86_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4267_ _0629_ _0939_ _0941_ mod.P3.Res\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_86_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6006_ _2535_ _2622_ _2624_ _2611_ _2625_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_80_1183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4198_ _0807_ mod.Arithmetic.CN.I_in\[26\] _0873_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_95_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_1219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_677 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_7957_ _0183_ net1 mod.Data_Mem.F_M.MRAM\[769\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1228 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1239 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6908_ _3379_ _0210_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4975__A1 mod.Data_Mem.F_M.MRAM\[6\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4913__S _1581_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_165_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7888_ _0114_ net1 mod.Data_Mem.F_M.MRAM\[25\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_23_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7213__I0 _3529_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6839_ _3246_ mod.Data_Mem.F_M.MRAM\[769\]\[3\] _3340_ _3342_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__4027__I0 _0638_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5924__B1 _2536_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8509_ net189 net1 mod.Data_Mem.F_M.out_data\[69\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__5029__B _1558_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3950__A2 mod.P2.Rout_reg\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5152__A1 _1574_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5455__A2 _2103_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5699__B _2259_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3998__I mod.Arithmetic.CN.I_in\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_611 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3120 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_19_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3131 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8506__D _0010_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3142 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3153 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_975 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6404__A1 _3009_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3164 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_85 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6404__B2 _2503_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3175 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2430 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3186 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2441 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3197 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2452 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2463 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2474 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4966__A1 _1620_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2485 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1740 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2496 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1751 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4966__B2 mod.Data_Mem.F_M.MRAM\[15\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1762 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1773 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1784 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_1795 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7755__I1 mod.Data_Mem.F_M.MRAM\[796\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_393 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6042__C _2659_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5391__A1 _1704_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4194__A2 _0804_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8532__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_465 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_128_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_115_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5453__I _2101_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5694__A2 _2140_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_714 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5170_ _1835_ _1836_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_69_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4121_ _0797_ _0747_ _0798_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_64_1167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_717 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4249__A3 _0660_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4052_ _0722_ _0721_ _0729_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_49_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_611 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_931 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xtiny_user_project_90 la_data_out[11] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_64_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_964 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_65_975 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7811_ mod.Data_Mem.F_M.MRAM\[7\]\[5\] _3904_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_64_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5829__S _2452_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7742_ mod.Data_Mem.F_M.MRAM\[795\]\[7\] _3865_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_52_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8062__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4957__A1 _1501_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4954_ _1620_ mod.Data_Mem.F_M.MRAM\[799\]\[0\] _1621_ mod.Data_Mem.F_M.MRAM\[783\]\[0\]
+ _1622_ _1623_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_33_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7673_ _3830_ _0524_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6233__B _2846_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4885_ mod.Data_Mem.F_M.src\[2\] _1554_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_71_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6624_ _3202_ _0103_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_20_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_933 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6555_ _3152_ _3153_ _3154_ _3155_ _3156_ _3157_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_69_1001 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_977 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_106_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5506_ _1677_ mod.Data_Mem.F_M.MRAM\[799\]\[6\] _2149_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_118_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4980__I1 mod.Data_Mem.F_M.MRAM\[2\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6486_ _3026_ _2309_ _3030_ _2497_ _2502_ _2672_ _3092_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_69_1056 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8225_ _0326_ net1 mod.Data_Mem.F_M.MRAM\[29\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_69_1078 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5437_ _2088_ _2089_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_160_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_1212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5685__A2 mod.Data_Mem.F_M.MRAM\[29\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5368_ _1888_ _2029_ _1863_ _2030_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_8156_ mod.Data_Mem.F_M.out_data\[66\] net2 net1 mod.Arithmetic.CN.I_in\[66\] vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_126_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7107_ _3500_ _3501_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_4319_ _0929_ _0658_ _0838_ _0993_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_101_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5299_ _1631_ _1949_ _1962_ _1963_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_8087_ _0287_ net1 mod.Data_Mem.F_M.MRAM\[23\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_75_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_47_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7038_ _3234_ _3464_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_47_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5312__B _1863_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8405__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_975 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6127__C _2743_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4660__A3 _1090_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_1016 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6398__B1 _3006_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6398__C2 _2510_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1014 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1025 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1036 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_35_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4948__A1 _1563_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5966__C _2263_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1058 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1069 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_168_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_42_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8555__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5538__I _2177_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_169_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_129_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_156_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_1082 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4176__A2 _0851_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5474__S _1908_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_1101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_87_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6322__B1 _2933_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_1178 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_809 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_319 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_980 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5920__I0 mod.Data_Mem.F_M.MRAM\[784\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_588 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_150_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_19_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4100__A2 _0773_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4617__I mod.Arithmetic.CN.I_in\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8085__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4651__A3 _1321_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_1149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2260 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_34_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2271 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2282 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2293 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5600__A2 _2221_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4403__A3 _0980_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_319 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1570 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1050 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_14_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1581 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5448__I _2096_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_159_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5739__I0 mod.Data_Mem.F_M.MRAM\[4\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4670_ _1339_ _1337_ _1340_ _1341_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__7922__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6561__B1 _3023_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6340_ _2886_ _2947_ _2950_ _2951_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_51_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6271_ _2837_ _2884_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_66_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8010_ _0219_ net1 mod.Data_Mem.F_M.MRAM\[14\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5222_ mod.Data_Mem.F_M.MRAM\[31\]\[4\] _1886_ _1887_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5153_ mod.Data_Mem.F_M.MRAM\[17\]\[3\] mod.Data_Mem.F_M.MRAM\[16\]\[3\] _1816_ _1819_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_96_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8428__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4104_ mod.Arithmetic.ACTI.x\[4\] _0781_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_84_503 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5419__A2 _2074_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5084_ _1524_ _1751_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_99_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4035_ _0684_ _0711_ _0702_ _0712_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__6092__A2 _1613_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4642__A3 mod.Arithmetic.CN.I_in\[30\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8578__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_169_107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_53_978 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_5986_ mod.Data_Mem.F_M.MRAM\[784\]\[5\] mod.Data_Mem.F_M.MRAM\[785\]\[5\] _1686_
+ _2606_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XPHY_119 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__7592__A2 _3446_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7725_ _3856_ _0550_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_40_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4937_ _1572_ _1606_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_36_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7774__S _3883_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7656_ mod.Data_Mem.F_M.MRAM\[790\]\[4\] _3822_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_138_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4868_ _1528_ _1537_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6607_ mod.Data_Mem.F_M.MRAM\[11\]\[7\] _3194_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5355__A1 _2012_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4158__A2 _0833_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_165_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_7587_ _3782_ mod.Data_Mem.F_M.MRAM\[785\]\[6\] _3779_ _3783_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__5294__S _1783_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4799_ _1314_ _1176_ _1310_ _1468_ _1469_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_107_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6538_ _2447_ _2337_ _2631_ _2642_ _3140_ _3141_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_118_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5107__A1 _1563_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_755 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_79 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6469_ _2151_ mod.Data_Mem.F_M.MRAM\[13\]\[3\] _3075_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_106_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_161_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_8208_ _0309_ net1 mod.Data_Mem.F_M.MRAM\[12\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_115_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8139_ mod.Data_Mem.F_M.out_data\[49\] net2 net1 mod.Arithmetic.CN.I_in\[49\] vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_43_1037 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_75_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_536 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_169_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4094__A1 _0747_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7945__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5594__A1 _2228_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4397__A2 mod.Arithmetic.CN.I_in\[28\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_169_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5268__I _1890_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_538 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4149__A2 mod.Arithmetic.CN.I_in\[48\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7483__I _3717_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5897__A2 _2509_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_939 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_125_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_606 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_617 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_639 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_152_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_1104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_864 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_1159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_856 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_93_344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_761 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5821__A2 _2444_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_539 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5379__S _1903_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_1093 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5840_ _2085_ _2446_ _2463_ _1498_ _0057_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_35_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_1200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_797 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2090 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5585__A1 _2221_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5771_ _2395_ _2396_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_99_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_61_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7594__S _3787_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7510_ _3735_ _0456_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4722_ _1269_ _1391_ _1393_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_8490_ _0586_ net1 mod.Data_Mem.F_M.MRAM\[7\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_33_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7441_ mod.Data_Mem.F_M.MRAM\[777\]\[5\] _3694_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_30_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8100__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5337__B2 _1999_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4653_ _1285_ _1323_ _1324_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_147_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5906__I _1894_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7372_ _3659_ _0394_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4935__I1 mod.Data_Mem.F_M.MRAM\[788\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4584_ _1236_ _1255_ _1256_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_128_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6230__C _2843_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6323_ _2920_ _2923_ _2930_ _2934_ _2935_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_116_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8250__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6254_ _2702_ _2867_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_5205_ mod.Data_Mem.F_M.MRAM\[15\]\[4\] _1870_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_130_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6185_ _1834_ _2799_ _2800_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5136_ _1695_ _1802_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_85_823 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_171 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7769__S _3878_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5067_ _1526_ _1734_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_38_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7968__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4018_ mod.Arithmetic.CN.I_in\[22\] _0695_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_65_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_25_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_285 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4379__A2 _0804_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5969_ _2588_ mod.Data_Mem.F_M.MRAM\[4\]\[5\] _2589_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_52_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7708_ mod.Data_Mem.F_M.MRAM\[793\]\[6\] _3848_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_32_23 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_139_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7317__A2 _3626_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7639_ _3813_ _0507_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_148_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7009__S _3440_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4551__A2 _1113_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6828__A1 mod.Data_Mem.F_M.dest\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_79_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_1159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4303__A2 _0933_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_121_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_983 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_171 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__6056__A2 _2673_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4067__A1 mod.Arithmetic.CN.I_in\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4067__B2 _0743_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_1192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_63_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_63_539 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8514__D _0018_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7556__A2 _3762_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_572 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8123__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5567__A1 mod.Data_Mem.F_M.MRAM\[29\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5567__B2 mod.Data_Mem.F_M.MRAM\[28\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5319__A1 _1551_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_1015 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_1086 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_117_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8273__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_156_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6119__I0 mod.Data_Mem.F_M.MRAM\[23\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4542__A2 mod.Arithmetic.CN.I_in\[36\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_101_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_469 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_121_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_536 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_27_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7990_ mod.Instr_Mem.instruction\[23\] net2 net1 mod.Data_Mem.F_M.src\[1\] vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_66_355 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6941_ _3253_ mod.Data_Mem.F_M.MRAM\[14\]\[5\] _3400_ _3402_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_66_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6292__I _1493_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6872_ _3358_ _0195_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_35_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5823_ _2352_ _2447_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5558__A1 _2189_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5558__B2 _1915_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8542_ _0046_ net1 mod.Data_Mem.F_M.out_data\[38\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5754_ _2378_ _2379_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4705_ _0632_ mod.Arithmetic.ACTI.x\[6\] _1376_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__6507__B1 _2500_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8473_ _0569_ net1 mod.Data_Mem.F_M.MRAM\[797\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5685_ _2313_ mod.Data_Mem.F_M.MRAM\[29\]\[4\] _2314_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__6507__C2 _2568_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6241__B _2733_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7424_ _3685_ _0420_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4636_ _1178_ _1307_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_118_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_7355_ mod.Data_Mem.F_M.MRAM\[772\]\[2\] _3651_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4567_ _1126_ _1130_ _1239_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_162_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6306_ _2876_ _1973_ _2763_ _2918_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_7286_ _3607_ _0360_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4696__B _1366_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4498_ _1069_ _1071_ _1068_ _1170_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_89_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6286__A2 _2896_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6237_ _1931_ _1848_ _2851_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_131_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5333__I1 mod.Data_Mem.F_M.MRAM\[18\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8527__179 net179 vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XANTENNA__4297__A1 _0618_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_801 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6168_ _2779_ _2780_ _2783_ _2692_ _2784_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_112_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_981 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7499__S _3726_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5119_ _1782_ mod.Data_Mem.F_M.MRAM\[789\]\[2\] _1785_ _1786_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_45_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6099_ _2195_ _2711_ _2712_ _2715_ _2716_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_17_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6443__C1 _2460_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2804 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2815 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_539 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5797__A1 _2110_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8146__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2826 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2837 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2848 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2859 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6210__A2 _1786_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8296__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4221__A1 _0643_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_1196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_166_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_138_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_154_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5721__A1 _2312_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4524__A2 _1187_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_122_500 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_136_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5324__I1 mod.Data_Mem.F_M.MRAM\[4\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_150_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_74 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_823 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_290 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5788__A1 _1490_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_1030 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_147_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4460__A1 _1124_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4212__A1 _0825_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_291 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__4763__A2 _1354_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5470_ _2117_ _2118_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_157_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_8_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8194__RN net2 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4421_ _1092_ _1093_ _1094_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__8019__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_99_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7140_ _3520_ _0301_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_154_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4352_ _0948_ _1025_ _1026_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_113_533 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7071_ _3482_ _0270_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4283_ _0875_ _0956_ _0957_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__4279__A1 _0687_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5476__B1 _2119_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6022_ _2587_ mod.Data_Mem.F_M.MRAM\[5\]\[6\] _2640_ _2091_ _2641_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_98_288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8169__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7112__S _3501_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_984 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7973_ _0199_ net1 mod.Data_Mem.F_M.MRAM\[6\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_54_325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6236__B _2738_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4535__I _1206_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6924_ _3235_ _3387_ _3389_ _3390_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_70_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6440__A2 _2451_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6855_ mod.Data_Mem.F_M.MRAM\[779\]\[3\] _3350_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_50_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7240__I1 mod.Data_Mem.F_M.MRAM\[30\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5806_ _2358_ mod.Data_Mem.F_M.MRAM\[789\]\[1\] _2430_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_23_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6786_ _3305_ _3306_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_3998_ mod.Arithmetic.CN.I_in\[15\] _0675_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_8525_ net181 net1 mod.Data_Mem.F_M.out_data\[53\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__4754__A2 _1423_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5737_ _2162_ _2362_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_148_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_8456_ _0552_ net1 mod.Data_Mem.F_M.MRAM\[795\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_135_113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_108_327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5668_ _2068_ _2298_ _2299_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_11_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7407_ mod.Data_Mem.F_M.MRAM\[775\]\[4\] _3677_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_136_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4619_ _0737_ mod.Arithmetic.CN.I_in\[13\] _1190_ _1290_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__7581__I _3772_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8387_ _0483_ net1 mod.Data_Mem.F_M.MRAM\[785\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5599_ _1574_ _2235_ _2236_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_2_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_150_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_163_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_117_894 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7338_ _3641_ _0378_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_46_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_89_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7269_ mod.Data_Mem.F_M.MRAM\[5\]\[2\] _3597_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_104_588 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_58_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6925__I _3390_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_995 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2601 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2612 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2623 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_166_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2634 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_166_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2645 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1900 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2656 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1911 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4442__A1 mod.Arithmetic.CN.I_in\[50\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2667 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1922 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1933 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2678 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2689 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1944 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1955 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5477__S _1510_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_391 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1966 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1977 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7231__I1 mod.Data_Mem.F_M.MRAM\[30\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6195__A1 _2759_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1988 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1999 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5242__I0 mod.Data_Mem.F_M.MRAM\[769\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_16_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_55_1091 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5942__A1 _2560_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5276__I _1573_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4745__A2 mod.Arithmetic.CN.I_in\[71\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_167_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_127_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_103_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_1056 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_1078 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8176__RN net2 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6498__A2 _2318_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_155_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_79_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__8311__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7298__I1 mod.Data_Mem.F_M.MRAM\[768\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_1040 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_536 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_1073 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xtiny_user_project_130 la_data_out[51] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_141 la_data_out[62] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_48_152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8461__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xtiny_user_project_152 wbs_dat_o[5] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_48_163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xtiny_user_project_163 wbs_dat_o[16] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_92_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xtiny_user_project_174 wbs_dat_o[27] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_63_122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8100__RN net2 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4970_ _1635_ _1637_ _1638_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_63_177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5481__I0 mod.Data_Mem.F_M.MRAM\[30\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4984__A2 _1648_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_840 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6640_ _3210_ _0111_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6186__A1 mod.Data_Mem.F_M.MRAM\[13\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_165_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6571_ mod.I_addr\[2\] _3171_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__5933__A1 _2434_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8310_ _0406_ net1 mod.Data_Mem.F_M.MRAM\[774\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5522_ _2161_ mod.Data_Mem.F_M.MRAM\[30\]\[0\] mod.Data_Mem.F_M.MRAM\[31\]\[0\] _2162_
+ _2163_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_118_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_1216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8241_ _0337_ net1 mod.Data_Mem.F_M.MRAM\[30\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__8167__RN net2 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5453_ _2101_ _2102_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5914__I _2394_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_319 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4404_ _1049_ _1075_ _1076_ _1077_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_114_820 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8172_ mod.P2.dest_reg\[2\] net2 net1 mod.Data_Mem.F_M.dest\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_5384_ _1872_ _2045_ _1884_ _2046_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_113_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7123_ _3510_ _0294_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4335_ mod.Arithmetic.CN.I_in\[64\] _0918_ mod.Arithmetic.ACTI.x\[1\] _0643_ _1009_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XFILLER_99_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_875 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_119_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7054_ _3460_ mod.Data_Mem.F_M.MRAM\[1\]\[6\] _3469_ _3474_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_87_748 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6110__A1 _2185_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4266_ _0768_ _0855_ _0857_ _0940_ _0627_ _0941_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_80_1151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6745__I _3273_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6005_ _2062_ mod.Data_Mem.F_M.MRAM\[772\]\[6\] _2623_ _2624_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_80_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_461 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4197_ mod.Arithmetic.CN.I_in\[24\] _0871_ _0808_ _0872_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or3_1
XFILLER_80_1195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7956_ _0182_ net1 mod.Data_Mem.F_M.MRAM\[769\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1207 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4424__A1 _0897_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1229 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6907_ _3243_ mod.Data_Mem.F_M.MRAM\[13\]\[2\] _3376_ _3379_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_70_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_1080 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7887_ _0113_ net1 mod.Data_Mem.F_M.MRAM\[25\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__4975__A2 _1640_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7213__I1 mod.Data_Mem.F_M.MRAM\[2\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6838_ _3341_ _0178_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6177__A1 _2199_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4027__I1 mod.Arithmetic.I_out\[72\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6769_ _3291_ _0159_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_155_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5924__B2 _2538_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_149_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_8508_ net190 net1 mod.Data_Mem.F_M.out_data\[68\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_40_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8334__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8439_ _0535_ net1 mod.Data_Mem.F_M.MRAM\[792\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__8158__RN net2 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_156_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_3_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_151_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_680 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5152__A2 _1817_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_1046 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8484__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_759 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_962 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_59_984 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4663__A1 mod.Arithmetic.CN.I_in\[38\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3110 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3121 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3132 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3143 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3154 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3165 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2420 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_34_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_45_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6404__A2 _2389_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2431 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_678 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3176 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3187 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2442 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5463__I0 mod.Data_Mem.F_M.MRAM\[30\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_3198 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2453 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2464 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2475 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1730 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2486 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_121_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4966__A2 _1632_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_1153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1752 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2497 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1763 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4903__I _1571_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_1017 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1774 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1066 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6168__A1 _2779_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1785 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5215__I0 mod.Data_Mem.F_M.MRAM\[3\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_1197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1796 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_147_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_1129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4718__A2 _1388_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5935__S _2301_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5391__A2 _2052_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_127_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8149__RN net2 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6340__A1 _2886_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4120_ mod.P2.Rout_reg\[0\] _0797_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_68_214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_151_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_110_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_110_355 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4051_ _0725_ _0727_ _0728_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_68_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xtiny_user_project_80 la_data_out[1] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_91 la_data_out[12] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
X_7810_ _3903_ _0588_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_64_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_773 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__8207__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4406__A1 _0813_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_149_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_52_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_1220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7741_ _3864_ _0558_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_80_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4953_ _1550_ _1622_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__4957__A2 _1553_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6514__B _2406_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_162_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7672_ mod.Data_Mem.F_M.MRAM\[791\]\[4\] _3830_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4884_ _1534_ _1553_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_20_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6623_ mod.Data_Mem.F_M.MRAM\[24\]\[7\] _3202_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__8357__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6954__I0 _3393_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6554_ _2548_ _2673_ _3156_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_119_945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_5505_ _2135_ mod.Data_Mem.F_M.MRAM\[30\]\[6\] _2147_ _2148_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_134_915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6485_ _2072_ _2509_ _3086_ _3090_ _3091_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_161_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_106_639 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8224_ _0325_ net1 mod.Data_Mem.F_M.MRAM\[29\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_133_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5436_ _2069_ _2088_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_133_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_126_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_8155_ mod.Data_Mem.F_M.out_data\[65\] net2 net1 mod.Arithmetic.CN.I_in\[65\] vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_5367_ _2024_ _2026_ _2027_ _2028_ _1881_ _1590_ _2029_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_120_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_102_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7106_ _3433_ _3272_ _3407_ _3500_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_87_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4318_ _0910_ _0991_ _0927_ _0933_ _0992_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_8086_ _0286_ net1 mod.Data_Mem.F_M.MRAM\[23\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5298_ _1633_ _1960_ _1961_ _1962_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_101_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7037_ _3463_ _0255_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__7831__A1 _0612_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4249_ _0619_ mod.Arithmetic.CN.I_in\[57\] _0660_ _0924_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_102_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4645__A1 _1061_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_16_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_43_604 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6398__A1 _3005_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1004 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7300__S _3608_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6398__B2 _2407_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1015 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1037 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_7939_ _0165_ net1 mod.Data_Mem.F_M.MRAM\[799\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_43_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4948__A2 _1605_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_169_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1048 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1059 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_1050 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_11_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_1072 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_167_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_1094 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_13_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_109_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7874__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7122__I0 _3460_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_1204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_751 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_678 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_773 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6389__A1 mod.Data_Mem.F_M.MRAM\[781\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6389__B2 mod.Data_Mem.F_M.MRAM\[780\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2250 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2261 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2272 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2283 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2294 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7189__I0 _3523_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1571 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1062 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6053__C _2263_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1582 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1593 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_119_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6561__A1 mod.Data_Mem.F_M.MRAM\[781\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6561__B2 mod.Data_Mem.F_M.MRAM\[769\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5464__I _1803_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_115_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_1208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6313__A1 _1826_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6270_ _1895_ _1893_ _1742_ _2883_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_44_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_5221_ _1672_ _1886_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_88_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_131_929 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_155_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_1022 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5152_ _1574_ _1817_ _1818_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_97_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4103_ _0725_ _0778_ _0779_ _0780_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XANTENNA__5419__A3 _2077_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5083_ mod.Data_Mem.F_M.MRAM\[22\]\[2\] _1749_ _1641_ _1750_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_84_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4627__A1 _1185_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_526 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6228__C _2841_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4034_ mod.Arithmetic.I_out\[73\] _0711_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_65_751 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_773 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7120__S _3506_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5985_ mod.Data_Mem.F_M.MRAM\[786\]\[5\] mod.Data_Mem.F_M.MRAM\[787\]\[5\] _1515_
+ _2605_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XPHY_109 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__5052__A1 _1700_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7724_ mod.Data_Mem.F_M.MRAM\[794\]\[6\] _3856_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4936_ mod.Data_Mem.F_M.MRAM\[790\]\[0\] _1601_ _1603_ _1604_ _1605_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_33_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_162_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_33_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_166_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7655_ _3821_ _0515_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_21_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4867_ _1535_ _1536_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6606_ _3193_ _0094_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_20_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7586_ _3318_ _3782_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5355__A2 _2015_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6552__A1 _2417_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4798_ _1314_ _1176_ _1310_ _1467_ _1468_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_119_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7897__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6537_ _2071_ _2210_ _2636_ _2698_ _3140_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_106_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7790__S _3889_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_959 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6304__A1 _1664_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6468_ _3017_ mod.Data_Mem.F_M.MRAM\[1\]\[3\] _3031_ _3073_ _3074_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_8207_ _0308_ net1 mod.Data_Mem.F_M.MRAM\[12\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5419_ _2072_ _2074_ _2077_ _0009_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_82_1010 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5902__I1 mod.Data_Mem.F_M.MRAM\[3\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6399_ _3004_ _3007_ _3008_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_121_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8138_ mod.Data_Mem.F_M.out_data\[48\] net2 net1 mod.Arithmetic.CN.I_in\[48\] vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_88_843 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_504 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8069_ _0278_ net1 mod.Data_Mem.F_M.MRAM\[21\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_101_152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__8522__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7030__S _3457_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5549__I _1790_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5043__A1 _1707_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8072__D mod.P3.Res\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_1161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_1156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_129_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6918__I0 _3259_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_169_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6543__A1 _3106_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_607 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8052__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4321__A3 mod.Arithmetic.CN.I_in\[51\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_113_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_38_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_751 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5282__A1 _1826_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5887__C _2508_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5459__I _2107_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6064__B _1535_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_607 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_1089 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2080 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_1212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5770_ _1595_ _1554_ _2395_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_2091 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_50_949 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_159_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4721_ _1269_ _1391_ _1392_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XTAP_1390 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_148_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6909__I0 _3246_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7440_ _3693_ _0428_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_30_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5337__A2 _1992_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4652_ _1286_ _1322_ _1323_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__7582__I0 _3778_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7371_ mod.Data_Mem.F_M.MRAM\[773\]\[2\] _3659_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_128_561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4583_ _1237_ _1254_ _1255_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_116_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6322_ _2895_ _2932_ _2933_ _2898_ _1866_ _2934_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_115_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7334__I0 _3638_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6298__B1 _2157_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6253_ _2374_ _2866_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_66_1049 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5204_ _1802_ _1803_ _1869_ _0003_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_112_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6184_ _2070_ mod.Data_Mem.F_M.MRAM\[14\]\[2\] mod.Data_Mem.F_M.MRAM\[15\]\[2\] _2203_
+ _2799_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_69_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8545__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5135_ _1729_ _1627_ _1760_ _1670_ _1801_ _0002_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_97_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_995 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5066_ mod.Data_Mem.F_M.MRAM\[6\]\[2\] _1601_ _1641_ _1733_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__4076__A2 _0751_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4017_ _0679_ mod.Arithmetic.I_out\[77\] _0689_ _0692_ _0693_ _0694_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_4
XFILLER_77_1112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4871__I1 mod.Data_Mem.F_M.MRAM\[4\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5025__A1 _1692_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_607 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_1178 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_77_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6773__A1 mod.Data_Mem.F_M.dest\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5968_ _1685_ _2588_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_40_426 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7707_ _3847_ _0541_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4919_ _1587_ _1588_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_5899_ mod.Data_Mem.F_M.MRAM\[4\]\[3\] mod.Data_Mem.F_M.MRAM\[5\]\[3\] mod.Data_Mem.F_M.MRAM\[20\]\[3\]
+ mod.Data_Mem.F_M.MRAM\[21\]\[3\] _1918_ _1756_ _2521_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_138_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6525__A1 _2558_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7638_ mod.Data_Mem.F_M.MRAM\[788\]\[3\] _3813_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_20_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_165_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_154_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_101_1110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7569_ _3292_ _3771_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_140_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_572 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_107_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8075__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_161_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6928__I _3239_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_164_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_533 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_88_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7912__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_1160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6461__B1 _2536_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_816 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_710 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_90_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_56_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_765 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5567__A2 _2200_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_1021 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7308__A3 _3446_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4911__I _1579_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_157_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8418__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_153_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8568__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_426 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_426 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_393 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_66_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_643 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_26_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5255__A1 _1906_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6940_ _3401_ _0220_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_47_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6871_ mod.Data_Mem.F_M.MRAM\[6\]\[3\] _3358_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6055__I0 mod.Data_Mem.F_M.MRAM\[2\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6204__B1 _1762_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5822_ _2416_ _2433_ _2445_ _2446_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_22_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5558__A2 mod.Data_Mem.F_M.MRAM\[799\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8541_ _0045_ net1 mod.Data_Mem.F_M.out_data\[37\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5753_ _2377_ _2378_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__8098__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4821__I _1489_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_1075 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4704_ _0641_ mod.Arithmetic.ACTI.x\[5\] _1125_ _1375_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_31_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6507__A1 _3049_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8472_ _0568_ net1 mod.Data_Mem.F_M.MRAM\[797\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_30_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5684_ _1691_ _2313_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__6507__B2 _2543_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_147_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_136_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7423_ mod.Data_Mem.F_M.MRAM\[776\]\[4\] _3685_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4635_ _1058_ _1304_ _1305_ _1306_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_159_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_159_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7354_ _3650_ _0385_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_116_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4566_ _0618_ mod.Arithmetic.CN.I_in\[68\] _1238_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_116_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6305_ _1655_ _1974_ _2917_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_143_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7285_ _3603_ mod.Data_Mem.F_M.MRAM\[768\]\[0\] _3606_ _3607_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_131_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4497_ _1053_ _1167_ _1168_ _1169_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_104_759 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6236_ _2845_ _2847_ _2738_ _2849_ _2850_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__7935__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4297__A2 mod.Arithmetic.CN.I_in\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5494__A1 _1677_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_1171 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6684__S _3237_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_48 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6167_ _2708_ _2781_ _2782_ _2783_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XTAP_971 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_982 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_1019 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5118_ _1783_ _1784_ _1785_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_73_805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6098_ _2714_ _2715_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_57_367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6443__B1 _3050_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6443__C2 _2496_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2805 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5049_ _1715_ _1716_ _1717_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_2816 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5797__A2 _2420_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2827 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2838 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2849 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_25_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_25_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_80_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_90_1153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4221__A2 mod.Arithmetic.CN.I_in\[42\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_1126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7546__I0 _3731_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3980__A1 _0655_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5721__A2 _2154_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4524__A3 _1195_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5562__I _1542_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_1200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5485__A1 _2129_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5237__A1 _1901_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4906__I _1574_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_646 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5938__S _2189_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4460__A2 _1132_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4842__S _1510_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8240__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_1086 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4212__A2 _0849_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5737__I _2162_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_270 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_13_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_292 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_129_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3971__A1 _0639_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8390__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4420_ _0828_ mod.Arithmetic.CN.I_in\[35\] _0826_ _0892_ _1093_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XANTENNA__7958__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4351_ _0951_ _0976_ _1024_ _1025_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_119_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_1177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_7070_ mod.Data_Mem.F_M.MRAM\[20\]\[6\] _3482_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_63_1019 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4282_ _0806_ mod.Arithmetic.CN.I_in\[19\] _0956_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_113_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4279__A2 _0804_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5476__A1 _2074_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6021_ _2345_ mod.Data_Mem.F_M.MRAM\[4\]\[6\] _2640_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__5476__B2 _2121_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8526__180 net180 vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_82_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7972_ _0198_ net1 mod.Data_Mem.F_M.MRAM\[6\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_54_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_646 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_540 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6923_ _3388_ _3389_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_165_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6854_ _3349_ _0186_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__7776__I0 _3806_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5805_ _2395_ _2429_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6785_ net5 _3305_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_3997_ mod.Arithmetic.CN.I_in\[23\] _0674_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_50_576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5251__I1 mod.Data_Mem.F_M.MRAM\[788\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_278 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5736_ mod.Data_Mem.F_M.MRAM\[16\]\[0\] mod.Data_Mem.F_M.MRAM\[17\]\[0\] _2360_ _2361_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_8524_ net182 net1 mod.Data_Mem.F_M.out_data\[52\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__7528__I0 _3718_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3962__A1 _0637_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8455_ _0551_ net1 mod.Data_Mem.F_M.MRAM\[794\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_108_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5667_ _2294_ _2296_ _2297_ _2298_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_164_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4618_ _1287_ _0724_ _1288_ _1289_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_7406_ _3676_ _0411_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_8386_ _0482_ net1 mod.Data_Mem.F_M.MRAM\[785\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5598_ _2233_ mod.Data_Mem.F_M.MRAM\[799\]\[4\] mod.Data_Mem.F_M.MRAM\[798\]\[4\]
+ _2234_ _2235_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
X_7337_ _3640_ mod.Data_Mem.F_M.MRAM\[771\]\[2\] _3636_ _3641_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4549_ _1122_ _1139_ _1221_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__5382__I _1607_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7268_ _3596_ _0353_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_104_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_131_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_89_256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8113__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_77_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6219_ _2567_ _2572_ mod.Data_Mem.F_M.MRAM\[20\]\[3\] _2833_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_7199_ _3533_ mod.Data_Mem.F_M.MRAM\[29\]\[4\] _3553_ _3557_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__7303__S _3608_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6427__B _2381_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_58_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6267__I0 _1889_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2602 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_890 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__8263__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2613 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2624 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2635 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_819 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1901 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2646 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2657 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1912 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4442__A2 _1114_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2668 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1923 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2679 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1934 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_584 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1945 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_159_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7767__I0 _3303_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1956 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1967 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1978 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1989 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5242__I1 mod.Data_Mem.F_M.MRAM\[768\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_166_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_127_615 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_142_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_154_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_5_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_122_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_716 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_80 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7213__S _3562_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xtiny_user_project_120 la_data_out[41] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_131 la_data_out[52] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_62_1085 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
Xtiny_user_project_142 la_data_out[63] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_64_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_985 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4681__A2 _0995_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xtiny_user_project_153 wbs_dat_o[6] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_97_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xtiny_user_project_164 wbs_dat_o[17] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_110_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtiny_user_project_175 wbs_dat_o[28] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_91_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6186__A2 _2200_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4197__A1 mod.Arithmetic.CN.I_in\[24\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6570_ _3170_ _0081_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5933__A2 _2553_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5521_ _1812_ _2162_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_160_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_74_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_121_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_157_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8240_ _0336_ net1 mod.Data_Mem.F_M.MRAM\[30\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5452_ _2008_ _1554_ _2101_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__5697__A1 _2256_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8136__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4403_ _0893_ _0829_ _0980_ _1076_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
X_8171_ mod.P2.dest_reg\[1\] net2 net1 mod.Data_Mem.F_M.dest\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_5383_ _2040_ _2041_ _2042_ _2043_ _2044_ _1590_ _2045_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_114_843 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_7122_ _3460_ mod.Data_Mem.F_M.MRAM\[3\]\[6\] _3506_ _3510_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__5135__C _1801_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4334_ _0640_ mod.Arithmetic.CN.I_in\[67\] _1008_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_99_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5449__A1 _1951_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7053_ _1971_ _3466_ _3473_ _0261_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_101_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4265_ _0768_ _0773_ _0794_ _0940_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_101_526 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8286__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6004_ _2588_ mod.Data_Mem.F_M.MRAM\[773\]\[6\] _2623_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__6247__B _2202_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4196_ mod.Arithmetic.CN.I_in\[26\] _0871_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_27_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7955_ _0181_ net1 mod.Data_Mem.F_M.MRAM\[769\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_43_819 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_70_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1208 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5621__A1 mod.Data_Mem.F_M.MRAM\[797\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1219 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5621__B2 mod.Data_Mem.F_M.MRAM\[796\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6906_ _3378_ _0209_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_7886_ _0112_ net1 mod.Data_Mem.F_M.MRAM\[25\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_126_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6837_ _3243_ mod.Data_Mem.F_M.MRAM\[769\]\[2\] _3340_ _3341_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_11_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6177__A2 _2682_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6768_ mod.Data_Mem.F_M.MRAM\[8\]\[7\] _3291_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_7_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5924__A2 _2140_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_148_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_8507_ _0011_ net1 mod.Data_Mem.F_M.out_data\[67\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5719_ _1714_ _2345_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6699_ _3248_ _3249_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_109_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8438_ _0534_ net1 mod.Data_Mem.F_M.MRAM\[792\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_136_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_607 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5688__A1 _2315_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_163_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_8369_ _0465_ net1 mod.Data_Mem.F_M.MRAM\[783\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_102_1090 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6001__I _1681_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4360__A1 _0780_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_160_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_104_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7033__S _3457_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4112__A1 _0743_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_93_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_59_974 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5860__A1 _2474_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3100 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8075__D mod.P3.Res\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3111 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3122 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3133 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3144 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3155 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2410 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3166 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2421 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3177 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2432 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3188 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2443 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8094__RN net2 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2454 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5463__I1 mod.Data_Mem.F_M.MRAM\[31\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3199 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8009__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1720 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2465 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2476 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1731 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2487 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1742 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2498 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1753 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_1764 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1775 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5287__I _1816_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_1029 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1786 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5215__I1 mod.Data_Mem.F_M.MRAM\[2\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1797 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8159__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_167_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_139_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_155_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5679__A1 _2089_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_29_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_64_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_868 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5151__I0 mod.Data_Mem.F_M.MRAM\[19\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4050_ _0726_ _0690_ _0713_ _0727_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_65_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xtiny_user_project_70 io_out[29] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_65_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtiny_user_project_81 la_data_out[2] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_83_229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xtiny_user_project_92 la_data_out[13] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_49_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_64_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_92_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5603__A1 _2228_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7740_ mod.Data_Mem.F_M.MRAM\[795\]\[6\] _3864_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4952_ _1507_ _1621_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_17_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7671_ _3829_ _0523_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5197__I _1557_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4883_ _1551_ _1552_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6622_ _3201_ _0102_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6954__I1 mod.Data_Mem.F_M.MRAM\[15\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6553_ _2343_ mod.Data_Mem.F_M.MRAM\[13\]\[7\] _2381_ _3155_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_5504_ _1791_ mod.Data_Mem.F_M.MRAM\[31\]\[6\] _2147_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_134_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6484_ _3030_ _2514_ _3089_ _3090_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_106_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8223_ _0324_ net1 mod.Data_Mem.F_M.MRAM\[29\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5435_ _2063_ _0010_ _0024_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_145_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_156_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_640 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4342__A1 _1007_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5366_ mod.Data_Mem.F_M.MRAM\[7\]\[7\] mod.Data_Mem.F_M.MRAM\[6\]\[7\] _1877_ _2028_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_8154_ mod.Data_Mem.F_M.out_data\[64\] net2 net1 mod.Arithmetic.CN.I_in\[64\] vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_99_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_99_362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7105_ _3499_ _0287_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4317_ _0921_ _0926_ _0991_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_99_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_59_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8085_ _0285_ net1 mod.Data_Mem.F_M.MRAM\[23\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_102_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5297_ mod.Data_Mem.F_M.MRAM\[783\]\[5\] _1599_ _1961_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_87_535 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6095__A1 _2196_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5142__I0 mod.Data_Mem.F_M.MRAM\[5\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7036_ _3462_ mod.Data_Mem.F_M.MRAM\[18\]\[7\] _3457_ _3463_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4248_ _0922_ _0923_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_68_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5842__A1 _2418_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7788__S _3889_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6692__S _3237_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_782 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4179_ _0854_ _0855_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_167_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8076__RN net2 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6398__A2 _2261_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_71_936 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1016 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_7938_ _0164_ net1 mod.Data_Mem.F_M.MRAM\[799\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_70_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1049 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_7869_ _0095_ net1 mod.Data_Mem.F_M.MRAM\[11\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__8301__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_169_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_168_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7028__S _3457_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8451__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_87_1158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6322__A2 _2932_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4333__A1 _0914_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_105_651 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7122__I1 mod.Data_Mem.F_M.MRAM\[3\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5503__C _2104_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_31 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7822__A2 _3169_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_730 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_1129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2240 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_34_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2251 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2262 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2273 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2284 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2295 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1550 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7189__I1 mod.Data_Mem.F_M.MRAM\[29\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1572 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_822 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_90 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1583 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1594 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__6546__C1 _2616_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_1151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_1162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6561__A2 _2596_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_1184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4572__A1 _0614_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_927 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_938 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_127_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_109_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6313__A2 _1952_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5220_ _1872_ _1883_ _1884_ _1885_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__4324__A1 _0930_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5372__I0 mod.Data_Mem.F_M.MRAM\[19\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4324__B2 _0997_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5151_ mod.Data_Mem.F_M.MRAM\[19\]\[3\] mod.Data_Mem.F_M.MRAM\[18\]\[3\] _1816_ _1817_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__6576__I _3174_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6077__A1 _2087_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4102_ _0727_ _0766_ _0779_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5082_ _1600_ _1749_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_57_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4627__A2 _1093_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4033_ _0709_ _0710_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__8324__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5984_ _2424_ mod.Data_Mem.F_M.MRAM\[789\]\[5\] _2603_ _2604_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_7723_ _3855_ _0549_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4935_ mod.Data_Mem.F_M.MRAM\[789\]\[0\] mod.Data_Mem.F_M.MRAM\[788\]\[0\] _1568_
+ _1604_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_36_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_1035 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7654_ mod.Data_Mem.F_M.MRAM\[790\]\[3\] _3821_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__8474__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4866_ _1534_ _1535_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6605_ mod.Data_Mem.F_M.MRAM\[11\]\[6\] _3193_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_7585_ _3781_ _0485_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6552__A2 mod.Data_Mem.F_M.MRAM\[12\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4012__B1 _0682_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4797_ _1312_ _1316_ _1467_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__8230__RN net2 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6536_ _2474_ _3134_ _3138_ _3139_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_118_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6467_ _2171_ mod.Data_Mem.F_M.MRAM\[0\]\[3\] _3073_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__6304__A2 _1970_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8206_ _0307_ net1 mod.Data_Mem.F_M.MRAM\[12\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5418_ _2076_ _2077_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6398_ _3005_ _2261_ _3006_ _2407_ _2404_ _2510_ _3007_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_115_971 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_1180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8137_ mod.Data_Mem.F_M.out_data\[47\] net2 net1 mod.Arithmetic.CN.I_in\[47\] vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_87_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5349_ _1602_ _2012_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_114_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6068__A1 _1676_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4079__B1 _0721_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8068_ _0277_ net1 mod.Data_Mem.F_M.MRAM\[21\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_82_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7019_ _3451_ _0249_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4935__S _1568_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_23 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_28_432 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6240__A1 _2160_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_169_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_54_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_788 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_169_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_1124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6918__I1 mod.Data_Mem.F_M.MRAM\[13\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_1168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_11_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6170__B _2739_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6543__A2 mod.Data_Mem.F_M.MRAM\[769\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_398 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_109_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_3_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4306__A1 _0891_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7991__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_127_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_152_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6396__I _2092_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8528__D _0032_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_844 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__8347__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5806__A1 _2358_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4609__A2 _1257_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7221__S _3567_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_432 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6345__B _2763_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_46_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_74_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7020__I _3242_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_1057 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8497__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_755 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6231__A1 _2169_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2070 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2081 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2092 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_62_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4720_ _1272_ _1390_ _1391_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__4793__A1 _1422_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1380 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1391 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6909__I1 mod.Data_Mem.F_M.MRAM\[13\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4651_ _1297_ _1300_ _1321_ _1322_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XANTENNA__4545__A1 _1213_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7370_ _3658_ _0393_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4582_ _1249_ _1253_ _1254_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_162_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6321_ _1943_ _1945_ _2044_ _2933_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_115_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6298__A1 mod.Data_Mem.F_M.MRAM\[781\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6252_ _2534_ _2844_ _2863_ _2865_ _0067_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_89_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_716 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_278 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5203_ _1631_ _1862_ _1868_ _1869_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_69_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6183_ _2206_ _2682_ _2798_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_97_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5134_ _1777_ _1798_ _1800_ _1801_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_97_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6845__I0 _3256_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_538 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5065_ _1730_ _1731_ _1732_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_84_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6470__A1 _2275_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4016_ _0690_ _0691_ _0693_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_37_251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_53_755 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6222__A1 _1734_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_574 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7864__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5967_ _2214_ _2587_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_80_596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7706_ mod.Data_Mem.F_M.MRAM\[793\]\[5\] _3847_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4784__A1 _0743_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4918_ _1586_ _1587_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_166_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5981__B1 _2600_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5898_ _2118_ _2505_ _2519_ _2520_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_7637_ _3812_ _0506_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6525__A2 _2598_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4849_ _1517_ _1518_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4536__A1 _0651_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7568_ _3770_ _0479_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_107_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6519_ _3120_ _3122_ _3123_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_146_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_7499_ _3645_ mod.Data_Mem.F_M.MRAM\[781\]\[5\] _3726_ _3728_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_106_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7306__S _3608_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_103_930 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5988__C _2607_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7041__S _3466_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6461__B2 _2486_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_169_1049 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_1_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_571 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7261__I0 mod.Data_Mem.F_M.MRAM\[31\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4775__A1 _1300_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_145_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_169_462 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_156_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_40_983 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4527__A1 _1108_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_144_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5327__I0 mod.Data_Mem.F_M.MRAM\[3\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_427 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_39_505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_1094 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_1037 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5255__A2 mod.Data_Mem.F_M.MRAM\[786\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6452__A1 _2345_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_94_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_93_165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7887__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_891 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_81_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6870_ _3357_ _0194_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_35_755 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6204__A1 _1566_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7252__I0 mod.Data_Mem.F_M.MRAM\[31\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6055__I1 mod.Data_Mem.F_M.MRAM\[3\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6204__B2 _1555_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5821_ _2434_ _2444_ _2445_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_50_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8540_ _0044_ net1 mod.Data_Mem.F_M.out_data\[36\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_50_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4766__A1 _1422_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5752_ _2106_ _2376_ _2377_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_148_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4703_ mod.Arithmetic.CN.I_in\[67\] _1245_ _0634_ mod.Arithmetic.ACTI.x\[4\] _1374_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
X_8471_ _0567_ net1 mod.Data_Mem.F_M.MRAM\[796\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_30_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6507__A2 _2323_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5683_ _2311_ _2312_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_124_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7422_ _3684_ _0419_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5715__B1 _2341_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4634_ _1170_ _1171_ _1180_ _1181_ _1305_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_163_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7353_ mod.Data_Mem.F_M.MRAM\[772\]\[1\] _3650_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5191__A1 _1836_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8512__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4565_ _1124_ _1132_ _1133_ _1138_ _1237_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_128_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6304_ _1664_ _1970_ _2873_ _2916_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__5318__I0 _1978_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_716 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7284_ _3605_ _3606_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_4496_ _1054_ _1056_ _1067_ _1072_ _1168_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_104_738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6235_ _2160_ _1827_ _2718_ _2848_ _2849_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_131_546 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5494__A2 mod.Data_Mem.F_M.MRAM\[799\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_950 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_83_1183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6166_ _1730_ _1711_ _2782_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_961 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_972 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_983 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_994 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5117_ mod.Data_Mem.F_M.MRAM\[788\]\[2\] _1784_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_6097_ _2713_ _2714_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_85_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6443__A1 _3049_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_677 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7491__I0 _3640_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5048_ mod.Data_Mem.F_M.MRAM\[768\]\[1\] _1716_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__6443__B2 _2453_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2806 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_84_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2817 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_150_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2828 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_66_891 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2839 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_168_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6999_ _3438_ _0242_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_80_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8042__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4757__A1 _1422_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_167_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_1143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5329__B _1863_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_1165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7546__I1 mod.Data_Mem.F_M.MRAM\[783\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_103_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_154_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5706__B1 _2333_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3980__A2 _0656_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8192__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5182__A1 _1845_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_153_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_1050 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7036__S _3457_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_150_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8078__D mod.P3.Res\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_1078 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_95_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_75_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5237__A2 _1699_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6434__A1 _2343_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7482__I0 _3620_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_603 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_17_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6037__I1 mod.Data_Mem.F_M.MRAM\[783\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_71_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_71_393 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6115__S _1707_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_157_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8535__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_145_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_67_1112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4350_ _0978_ _0990_ _1023_ _1024_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_119_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_125_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4281_ _0877_ _0954_ _0955_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_67_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5476__A2 _2118_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6020_ _2185_ _2148_ _2638_ _2263_ _2639_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_79_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6425__A1 _3020_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7473__I0 _3711_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7971_ _0197_ net1 mod.Data_Mem.F_M.MRAM\[6\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_67_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8065__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6922_ mod.Data_Mem.F_M.dest\[1\] _3333_ _3388_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_54_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_390 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7225__I0 _3539_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6853_ mod.Data_Mem.F_M.MRAM\[779\]\[2\] _3349_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_62_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_680 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5928__I _2144_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6025__S _2360_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5804_ _1903_ _2428_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4739__A1 _1334_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6784_ _3304_ _0161_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_149_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3996_ mod.Arithmetic.ACTI.x\[7\] _0673_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_8523_ _0027_ net1 mod.Data_Mem.F_M.out_data\[51\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5735_ _1677_ _2360_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_50_588 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5864__S _2452_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7528__I1 mod.Data_Mem.F_M.MRAM\[783\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_8454_ _0550_ net1 mod.Data_Mem.F_M.MRAM\[794\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__3962__A2 mod.Arithmetic.CN.I_in\[24\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7902__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5666_ _2290_ _2124_ _2297_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_7405_ mod.Data_Mem.F_M.MRAM\[775\]\[3\] _3676_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4617_ mod.Arithmetic.CN.I_in\[14\] _1288_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_8385_ _0481_ net1 mod.Data_Mem.F_M.MRAM\[785\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5597_ _1811_ _2234_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_135_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_1212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7336_ _3305_ _3640_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4548_ _1122_ _1139_ _1220_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_7267_ mod.Data_Mem.F_M.MRAM\[5\]\[1\] _3596_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_81_1109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4479_ _1044_ _1045_ _1143_ _1151_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_89_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5467__A2 _2099_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_104_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6218_ _2212_ _2219_ _2508_ _2832_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_58_611 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7198_ _2213_ _3550_ _3556_ _0323_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_131_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6149_ _2706_ _2765_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8408__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6416__A1 _3014_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_752 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6267__I1 _1891_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_603 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2603 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2614 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2625 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2636 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_23 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2647 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1902 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2658 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1913 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2669 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_714 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1924 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8558__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1935 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1946 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_41_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1957 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_533 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1968 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_80_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1979 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5059__B _1726_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_1093 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_155_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_16_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5155__A1 _1557_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5573__I _2210_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4902__A1 _1528_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_69_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_49_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4917__I _1578_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_942 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xtiny_user_project_110 la_data_out[31] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XANTENNA__8088__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xtiny_user_project_121 la_data_out[42] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_48_132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xtiny_user_project_132 la_data_out[53] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XANTENNA__6407__A1 _3003_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xtiny_user_project_143 user_irq[0] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_76_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtiny_user_project_154 wbs_dat_o[7] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_76_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xtiny_user_project_165 wbs_dat_o[18] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_64_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_1127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xtiny_user_project_176 wbs_dat_o[29] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_149_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_149_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5091__B1 _1721_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7925__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_588 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_897 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4197__A2 _0871_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5394__A1 mod.Data_Mem.F_M.MRAM\[799\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_1182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5520_ _1942_ _2161_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_8_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_67_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5451_ _1535_ _2100_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_117_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5483__I _2096_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5697__A2 mod.Data_Mem.F_M.MRAM\[29\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4402_ _1052_ _1074_ _1075_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_8170_ mod.P2.dest_reg\[0\] net2 net1 mod.Data_Mem.F_M.dest\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_5382_ _1607_ _2044_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__4099__I _0775_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7121_ _3509_ _0293_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_99_533 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4333_ _0914_ _1005_ _1006_ _1007_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_141_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_125_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7052_ _3316_ _3466_ _3473_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_4264_ _0861_ _0938_ _0939_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_87_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_588 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6110__A3 _2726_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6003_ _2619_ mod.Data_Mem.F_M.MRAM\[782\]\[6\] _2621_ _2622_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_68_942 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4121__A2 _0747_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4195_ _0638_ _0805_ _0869_ _0810_ _0870_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_67_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6247__C _2210_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_67_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7954_ _0180_ net1 mod.Data_Mem.F_M.MRAM\[769\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6905_ _3240_ mod.Data_Mem.F_M.MRAM\[13\]\[1\] _3376_ _3378_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_7885_ _0111_ net1 mod.Data_Mem.F_M.MRAM\[26\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_51_820 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6836_ _3336_ _3340_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_50_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_51_864 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_168_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4188__A2 _0822_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6767_ _3290_ _0158_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_3979_ mod.Arithmetic.CN.I_in\[40\] _0656_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_13_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8506_ _0010_ net1 mod.Data_Mem.F_M.out_data\[66\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_13_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5718_ _2343_ mod.Data_Mem.F_M.MRAM\[29\]\[7\] _2344_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_137_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6698_ net7 _3248_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5137__A1 _1669_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_164_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8437_ _0533_ net1 mod.Data_Mem.F_M.MRAM\[792\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5649_ _2060_ _2281_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_124_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5688__A2 mod.Data_Mem.F_M.MRAM\[28\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_8368_ _0464_ net1 mod.Data_Mem.F_M.MRAM\[783\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_2_426 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_844 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_104_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7319_ _1851_ _3626_ _3629_ _0371_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_46_1015 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8299_ _0395_ net1 mod.Data_Mem.F_M.MRAM\[773\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_78_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8230__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_104_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_901 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3101 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3112 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_105_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_58_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3123 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8380__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3134 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3145 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2400 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3156 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2411 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2422 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3167 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7948__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3178 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2433 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3189 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2444 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5612__A2 mod.Data_Mem.F_M.MRAM\[799\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2455 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1710 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2466 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1721 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2477 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1732 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1743 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2488 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2499 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1754 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1765 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_875 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1776 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1787 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1798 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5679__A2 _2131_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_155_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_64_1104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_123_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_64_1137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_150_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_1159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_96_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7023__I _3245_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_569 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5151__I1 mod.Data_Mem.F_M.MRAM\[18\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xtiny_user_project_60 io_out[11] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_7_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtiny_user_project_71 io_out[30] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_37_603 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xtiny_user_project_82 la_data_out[3] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_77_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtiny_user_project_93 la_data_out[14] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_77_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7053__A1 _1971_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_40_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_617 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4406__A3 _0715_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_51_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_639 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4951_ _1619_ _1620_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_45_680 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_output3_I net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7670_ mod.Data_Mem.F_M.MRAM\[791\]\[3\] _3829_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4882_ _1550_ _1551_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_71_1108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6621_ mod.Data_Mem.F_M.MRAM\[24\]\[6\] _3201_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_33_897 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_123_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8103__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6564__B1 _2656_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6552_ _2417_ mod.Data_Mem.F_M.MRAM\[12\]\[7\] _3154_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_9_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_5503_ _2085_ _2142_ _2146_ _2104_ _0037_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XANTENNA__5119__A1 _1782_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6483_ _2439_ _3087_ _3088_ _3089_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XANTENNA__8253__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8222_ _0323_ net1 mod.Data_Mem.F_M.MRAM\[29\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5434_ _2080_ _2077_ _0019_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_127_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8153_ mod.Data_Mem.F_M.out_data\[63\] net2 net1 mod.Arithmetic.CN.I_in\[63\] vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_82_1204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4342__A2 _1015_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5390__I1 mod.Data_Mem.F_M.MRAM\[784\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5365_ mod.Data_Mem.F_M.MRAM\[5\]\[7\] mod.Data_Mem.F_M.MRAM\[4\]\[7\] _1877_ _2027_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__7134__S _3513_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7104_ mod.Data_Mem.F_M.MRAM\[23\]\[7\] _3499_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_87_503 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4316_ _0988_ _0989_ _0990_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_8084_ _0284_ net1 mod.Data_Mem.F_M.MRAM\[23\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5296_ _1622_ _1959_ _1960_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_7035_ _3258_ _3462_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_87_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5142__I1 mod.Data_Mem.F_M.MRAM\[4\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4247_ mod.Arithmetic.CN.I_in\[58\] _0922_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_101_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_68_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5842__A2 mod.Data_Mem.F_M.MRAM\[787\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4178_ _0672_ _0673_ _0854_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_68_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1006 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_83_797 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1017 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7937_ _0163_ net1 mod.Data_Mem.F_M.MRAM\[799\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_55_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7868_ _0094_ net1 mod.Data_Mem.F_M.MRAM\[11\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_169_836 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_169_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6819_ _3328_ _0172_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_7799_ _3322_ mod.Data_Mem.F_M.MRAM\[798\]\[7\] _3894_ _3898_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_7_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6440__C _3047_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_109_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_1126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5905__I0 mod.Data_Mem.F_M.MRAM\[14\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_152_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_105_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5851__I _1535_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_151_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7283__A1 _3232_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6330__I0 _2240_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_1181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_539 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_111_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2230 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2241 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__8126__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2252 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2263 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2274 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2285 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1540 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2296 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1551 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1562 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_80 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_14_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1573 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_91 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1584 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6546__B1 _2500_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1595 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_159_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6546__C2 _2568_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8276__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_128_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_755 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_1196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4572__A2 mod.Arithmetic.ACTI.x\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_155_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4324__A2 _0995_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5372__I1 mod.Data_Mem.F_M.MRAM\[18\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_503 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_111_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5150_ _1586_ _1816_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_96_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_151_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_611 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_536 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6078__B _1726_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4101_ _0746_ _0778_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_5081_ _1745_ _1747_ _1562_ _1748_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__4088__A1 _0748_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_355 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4032_ mod.Arithmetic.CN.I_in\[9\] _0709_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_38_923 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_24_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_797 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5588__A1 _1800_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5983_ _2398_ _1934_ _2603_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_64_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7722_ mod.Data_Mem.F_M.MRAM\[794\]\[5\] _3855_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_52_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4934_ _1602_ _1603_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5001__I mod.Data_Mem.F_M.src\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7329__A2 _3296_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7653_ _3820_ _0514_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4865_ mod.Data_Mem.F_M.src\[4\] _1534_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_6604_ _3192_ _0093_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_162_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7584_ _3754_ mod.Data_Mem.F_M.MRAM\[785\]\[5\] _3779_ _3781_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__4012__A1 _0680_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4012__B2 _0683_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4796_ _1302_ _1320_ _1465_ _1466_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_119_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6968__S _3414_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6535_ _3060_ _2643_ _2644_ _3020_ _3137_ _3138_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_118_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6466_ _3063_ _3072_ _0074_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_118_287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_427 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_133_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8205_ _0306_ net1 mod.Data_Mem.F_M.MRAM\[12\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__5512__A1 _2151_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5417_ _2075_ _2076_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_47_1110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5671__I _1692_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6397_ _2429_ _3006_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_86_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_983 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_114_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8136_ mod.Data_Mem.F_M.out_data\[46\] net2 net1 mod.Arithmetic.CN.I_in\[46\] vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_86_1192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5348_ _1700_ _2010_ _2011_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_749 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_87_322 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6068__A2 _2375_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8067_ _0276_ net1 mod.Data_Mem.F_M.MRAM\[21\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_102_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5279_ mod.Data_Mem.F_M.MRAM\[787\]\[5\] mod.Data_Mem.F_M.MRAM\[786\]\[5\] _1942_
+ _1943_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__4079__A1 _0754_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7018_ _3450_ mod.Data_Mem.F_M.MRAM\[18\]\[1\] _3448_ _3451_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_101_165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8149__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_83_572 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_797 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_70_233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6007__I _1757_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6240__A2 _1853_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8299__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4251__A1 _0923_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_24_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_1136 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_169_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_168_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4554__A2 _0995_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5782__S _1769_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_532 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5503__A1 _2085_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4306__A2 mod.Arithmetic.CN.I_in\[35\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_972 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_609 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_105_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_133_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7502__S _3726_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_1052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_19_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6231__A2 _1837_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2060 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_146_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2071 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_62_789 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4242__A1 _0615_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2082 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2093 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_981 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1370 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1381 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4793__A2 _1462_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5990__A1 _2079_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1392 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_642 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4650_ _1302_ _1320_ _1321_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_128_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4581_ _1018_ _1250_ _1136_ _1252_ _1253_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
X_6320_ _1566_ _1936_ _2931_ _2932_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_128_596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_157_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6298__A2 _2751_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6251_ _2079_ _2864_ _2865_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_88_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5202_ _1864_ _1865_ _1867_ _1699_ _1868_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_6182_ _2073_ _2792_ _2796_ _2797_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_130_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_69_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5133_ _1799_ _1800_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_112_964 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_675 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6845__I1 mod.Data_Mem.F_M.MRAM\[769\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5064_ mod.Data_Mem.F_M.MRAM\[5\]\[2\] mod.Data_Mem.F_M.MRAM\[4\]\[2\] _1636_ _1731_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_111_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4015_ _0690_ _0691_ _0680_ _0681_ _0692_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XFILLER_42_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8441__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5867__S _2452_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6222__A2 _1819_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5966_ _2579_ _2584_ _2585_ _2263_ _2586_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__4233__A1 _0662_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_52_277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7705_ _3846_ _0540_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4917_ _1578_ _1586_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5981__A1 _2596_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8591__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5981__B2 _2397_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5897_ _2416_ _2509_ _2518_ _2519_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_7636_ mod.Data_Mem.F_M.MRAM\[788\]\[2\] _3812_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_32_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4848_ _1512_ _1517_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_148_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_166_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7567_ _3731_ mod.Data_Mem.F_M.MRAM\[784\]\[7\] _3759_ _3770_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__4536__A2 mod.Arithmetic.CN.I_in\[45\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4779_ _1306_ _1318_ _1449_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_113_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6518_ _3111_ _3121_ _3122_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_101_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7498_ _3727_ _0452_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6449_ _3017_ mod.Data_Mem.F_M.MRAM\[781\]\[2\] _3056_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_162_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_103_942 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8119_ mod.Data_Mem.F_M.out_data\[29\] net2 net1 mod.Arithmetic.CN.I_in\[29\] vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_0_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7322__S _3625_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4847__I0 mod.Data_Mem.F_M.MRAM\[19\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_169_1017 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__6461__A2 _1886_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_1184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_84_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6960__I _3408_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7261__I1 _3319_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_789 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_575 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_1080 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4775__A2 _1321_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_995 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5724__A1 _2280_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4527__A2 _1140_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_1029 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__8314__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5327__I1 mod.Data_Mem.F_M.MRAM\[2\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5488__B1 _2131_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_152_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_1062 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__8464__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5335__S0 _1844_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_66_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5260__B _1674_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8130__RN net2 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6452__A2 _1770_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4463__A1 _0642_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_93_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6204__A2 _1761_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7252__I1 _3306_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5820_ _2435_ _2437_ _2438_ _2439_ _2443_ _2444_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_23_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4215__A1 _0830_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_1000 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5751_ _2375_ _2376_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_76_1191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5963__A1 _2397_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4766__A2 mod.Arithmetic.ACTI.x\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4390__I _1062_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4702_ _0643_ mod.Arithmetic.CN.I_in\[70\] _1373_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_8470_ _0566_ net1 mod.Data_Mem.F_M.MRAM\[796\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5682_ _2069_ _2311_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_7421_ mod.Data_Mem.F_M.MRAM\[776\]\[3\] _3684_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_148_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8197__RN net2 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5715__A1 _2082_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4633_ _1180_ _1181_ _1170_ _1171_ _1304_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XANTENNA__5715__B2 _2306_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_162_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7352_ _3649_ _0384_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5191__A2 mod.Data_Mem.F_M.MRAM\[769\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4564_ _1234_ _1235_ _1236_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_6303_ _2870_ _1969_ _2915_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_7283_ _3232_ _3332_ _3604_ _3605_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__5318__I1 _1979_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4495_ _1067_ _1072_ _1054_ _1056_ _1167_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_144_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5479__B1 _2125_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6234_ _2723_ _1830_ _2848_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__6140__A1 _2750_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_83_1151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6165_ _1706_ _1718_ _2781_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_951 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_962 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_69_152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_1195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_995 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5116_ _1567_ _1783_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_85_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_984 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_995 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6096_ _1500_ _1541_ _2713_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_131_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_57_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8121__RN net2 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6443__A2 _2285_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5047_ _1646_ _1715_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_2807 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_66_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4454__A1 _0915_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2818 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2829 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_84_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_81_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6998_ _3395_ mod.Data_Mem.F_M.MRAM\[17\]\[2\] _3435_ _3438_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__7981__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_13_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_748 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5949_ _2567_ mod.Data_Mem.F_M.MRAM\[2\]\[4\] _2568_ _2569_ _2570_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__5954__A1 _2506_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_1106 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_1188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8337__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_167_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5706__A1 _2082_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7619_ _3802_ _0498_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5706__B2 _2306_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5182__A2 mod.Data_Mem.F_M.MRAM\[773\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7116__I _3500_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8487__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6131__A1 _2169_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_569 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6682__A2 _3232_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_150_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_103_761 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_88_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_49_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_859 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6176__B _2791_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6434__A2 mod.Data_Mem.F_M.MRAM\[12\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7482__I1 mod.Data_Mem.F_M.MRAM\[780\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8112__RN net2 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_678 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6690__I net5 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_90_158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_1017 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_726 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5945__A1 _1533_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_31_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_9_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_169_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_76_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_144_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4220__I1 _0893_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_875 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_748 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_536 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4280_ _0871_ _0646_ _0809_ _0954_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_98_225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_98_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6865__I mod.Data_Mem.F_M.MRAM\[6\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4684__A1 mod.Arithmetic.CN.I_in\[52\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8103__RN net2 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7970_ _0196_ net1 mod.Data_Mem.F_M.MRAM\[6\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__4436__A1 _0930_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4436__B2 _0997_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6921_ _3373_ _3387_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_48_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7225__I1 mod.Data_Mem.F_M.MRAM\[2\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_165_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6852_ _3348_ _0185_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6189__A1 _2360_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6189__B2 _2188_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_1117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5803_ _2424_ _1678_ _2426_ _2427_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_90_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5936__A1 _2366_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6783_ mod.Data_Mem.F_M.MRAM\[799\]\[1\] _3303_ _3300_ _3304_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_167_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3995_ mod.P2.Rout_reg\[1\] _0672_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_22_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8522_ _0026_ net1 mod.Data_Mem.F_M.out_data\[50\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5734_ mod.Data_Mem.F_M.MRAM\[14\]\[0\] mod.Data_Mem.F_M.MRAM\[15\]\[0\] _2358_ _2359_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_8453_ _0549_ net1 mod.Data_Mem.F_M.MRAM\[794\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_149_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5665_ _2295_ mod.Data_Mem.F_M.MRAM\[28\]\[2\] _2259_ _2296_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__3962__A3 _0638_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7404_ _3675_ _0410_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_163_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_820 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4616_ mod.Arithmetic.CN.I_in\[13\] _1287_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_8384_ _0480_ net1 mod.Data_Mem.F_M.MRAM\[785\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5596_ _1594_ _2233_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5165__B _1614_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7335_ _3639_ _0377_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6976__S _3423_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4547_ _1205_ _1218_ _1219_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__5880__S _2339_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_150_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_117_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_104_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7266_ _3595_ _0352_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6113__A1 _2728_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_322 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7161__I0 _3533_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4478_ _1044_ _1045_ _1143_ _1150_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XANTENNA__7861__A1 _3917_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6217_ _2107_ _2831_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_132_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7197_ _3555_ _3550_ _3556_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_98_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6148_ _1640_ _2760_ _2762_ _2763_ _2764_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XTAP_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_781 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_645 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6079_ _2295_ _2696_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_100_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4427__A1 _1097_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2604 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2615 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2626 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2637 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2648 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1903 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2659 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1914 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1925 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_501 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1936 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1947 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_159_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1081 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1958 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1969 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_1092 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_41_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_70_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_103_1048 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7877__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4902__A2 _1541_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6104__A1 _2718_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4115__B1 _0789_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4666__A1 _1251_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_539 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_1054 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xtiny_user_project_100 la_data_out[21] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_0_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xtiny_user_project_111 la_data_out[32] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_88_291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xtiny_user_project_122 la_data_out[43] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_77_965 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xtiny_user_project_133 la_data_out[54] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_48_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xtiny_user_project_144 user_irq[1] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_155 wbs_dat_o[8] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XANTENNA__4418__A1 _0655_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xtiny_user_project_166 wbs_dat_o[19] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XANTENNA__5615__B1 _2249_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtiny_user_project_177 wbs_dat_o[30] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_76_497 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_92_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5091__A1 _1757_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8502__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5091__B2 mod.Data_Mem.F_M.MRAM\[15\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4933__I _1525_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_832 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6966__I0 _3403_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_149_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4197__A3 _0808_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_1194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5450_ _2097_ mod.Data_Mem.F_M.MRAM\[798\]\[0\] _2098_ _2099_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_161_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4401_ _1053_ _1057_ _1073_ _1074_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
X_5381_ mod.Data_Mem.F_M.MRAM\[775\]\[7\] mod.Data_Mem.F_M.MRAM\[774\]\[7\] _1908_
+ _2043_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_132_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_7120_ _3508_ mod.Data_Mem.F_M.MRAM\[3\]\[5\] _3506_ _3509_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4332_ _0665_ _0846_ _0919_ _1006_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or3_1
XANTENNA__7143__I0 _3462_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_99_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4106__B1 _0780_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7051_ _3472_ _0260_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5713__B _2311_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_4263_ _0862_ _0937_ _0938_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__8032__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4657__A1 _1206_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6002_ _2620_ mod.Data_Mem.F_M.MRAM\[783\]\[6\] _2621_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__6528__C _2079_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4194_ _0644_ _0804_ _0869_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_67_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_28_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_41_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_80_1187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7953_ _0179_ net1 mod.Data_Mem.F_M.MRAM\[769\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__8182__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_136 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_968 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6544__B _2474_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6904_ _3377_ _0208_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_7884_ _0110_ net1 mod.Data_Mem.F_M.MRAM\[26\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_63_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_1094 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_165_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_51_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6835_ _3339_ _0177_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_50_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5875__S _1932_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6766_ mod.Data_Mem.F_M.MRAM\[8\]\[6\] _3290_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4188__A3 _0669_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3978_ _0654_ _0655_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_50_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5717_ _1691_ _2343_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_8505_ _0009_ net1 mod.Data_Mem.F_M.out_data\[65\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_109_606 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6709__I0 _3256_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6697_ _3247_ _0131_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_108_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8436_ _0532_ net1 mod.Data_Mem.F_M.MRAM\[792\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_40_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5648_ _2088_ _2280_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6334__A1 _2870_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_156_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_8367_ _0463_ net1 mod.Data_Mem.F_M.MRAM\[782\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5579_ _2216_ _2217_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_151_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_2_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7318_ _3555_ _3623_ _3629_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__7134__I0 _3454_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8298_ _0394_ net1 mod.Data_Mem.F_M.MRAM\[773\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_2_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_104_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_46_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7249_ _3586_ _0344_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_86_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8525__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3102 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_615 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_784 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3113 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3124 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3135 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3146 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2401 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3157 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2412 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5073__A1 _1738_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3168 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2423 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3179 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2434 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4753__I mod.Arithmetic.CN.I_in\[38\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2445 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1700 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_164_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_73_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1711 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2456 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_1123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2467 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1722 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6173__C _2750_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2478 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1733 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2489 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_121_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_14_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1744 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1755 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1766 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1777 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1788 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1799 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_10_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_155_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_128_926 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_127_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__8055__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7505__S _3726_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4887__A1 _1553_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4351__A3 _1024_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_1127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4639__A1 _0844_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_526 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xtiny_user_project_50 io_out[1] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_61 io_out[12] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_72 io_out[31] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_49_464 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_76_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtiny_user_project_83 la_data_out[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_94 la_data_out[15] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XANTENNA__7240__S _3579_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7053__A2 _3466_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4950_ _1499_ _1619_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_17_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4406__A4 mod.Arithmetic.CN.I_in\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_1201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_938 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_1212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2990 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_36_1207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6939__I0 _3399_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4881_ _1548_ _1549_ _1550_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6620_ _3200_ _0101_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_60_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6564__A1 _2503_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6564__B2 _3050_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6551_ _2511_ mod.Data_Mem.F_M.MRAM\[0\]\[7\] _2103_ _3153_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_119_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5502_ _2143_ _2145_ _2084_ _2146_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__6316__A1 _2891_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6482_ _2475_ mod.Data_Mem.F_M.MRAM\[780\]\[3\] _3088_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_8221_ _0322_ net1 mod.Data_Mem.F_M.MRAM\[29\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_69_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5433_ _2085_ _2087_ _2076_ _0018_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_133_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4878__A1 _1508_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8152_ mod.Data_Mem.F_M.out_data\[62\] net2 net1 mod.Arithmetic.CN.I_in\[62\] vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_5364_ mod.Data_Mem.F_M.MRAM\[3\]\[7\] mod.Data_Mem.F_M.MRAM\[2\]\[7\] _2025_ _2026_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_160_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_1216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8548__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7103_ _3498_ _0286_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4315_ _0979_ _0987_ _0989_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_102_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8083_ _0283_ net1 mod.Data_Mem.F_M.MRAM\[23\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_113_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5295_ _1950_ _1952_ _1957_ _1958_ _1745_ _1822_ _1959_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_87_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7034_ _3461_ _0254_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_101_325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4246_ _0913_ _0920_ _0921_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_68_751 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4177_ _0801_ _0852_ _0853_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_95_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_67_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5055__A1 mod.Data_Mem.F_M.MRAM\[783\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6252__B1 _2863_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1007 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7936_ _0162_ net1 mod.Data_Mem.F_M.MRAM\[799\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1018 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1029 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_23_320 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7867_ _0093_ net1 mod.Data_Mem.F_M.MRAM\[11\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_168_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_23_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_504 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6818_ mod.Data_Mem.F_M.MRAM\[789\]\[4\] _3328_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_7798_ _3897_ _0582_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_50_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6749_ _3281_ _0149_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_137_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_109_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8078__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_1086 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4581__A3 _1136_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4318__B1 _0927_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8419_ _0515_ net1 mod.Data_Mem.F_M.MRAM\[790\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_87_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5905__I1 mod.Data_Mem.F_M.MRAM\[15\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6168__C _2692_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7915__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6330__I1 _2243_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_47_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6963__I _3252_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_773 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_1193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_968 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5579__I _2216_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2220 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_62_927 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2231 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2242 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2253 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2264 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1530 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2275 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2286 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1541 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2297 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1552 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_1032 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1563 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_81 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_30_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1574 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_92 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1585 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6546__A1 _3049_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6546__B2 _2615_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7594__I0 _3771_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_127_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7235__S _3574_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4100_ _0772_ _0773_ _0774_ _0776_ _0777_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_123_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5080_ mod.Data_Mem.F_M.MRAM\[19\]\[2\] mod.Data_Mem.F_M.MRAM\[18\]\[2\] _1746_ _1747_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_84_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4031_ _0682_ mod.Arithmetic.I_out\[74\] _0703_ _0708_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_96_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5489__I _2059_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_607 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5982_ mod.Data_Mem.F_M.MRAM\[770\]\[5\] mod.Data_Mem.F_M.MRAM\[771\]\[5\] _2522_
+ _2602_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_64_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_724 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_584 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_426 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7721_ _3854_ _0548_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4933_ _1525_ _1602_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_80_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_166_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7329__A3 _3634_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8220__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_1037 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6537__A1 _2071_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7652_ mod.Data_Mem.F_M.MRAM\[790\]\[2\] _3820_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4864_ _1496_ _1533_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_32_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_166_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_20_323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6603_ mod.Data_Mem.F_M.MRAM\[11\]\[5\] _3192_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_20_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7583_ _3780_ _0484_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_119_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4795_ _1303_ _1319_ _1465_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_6534_ _3135_ _3136_ _3137_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_146_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5157__C _1822_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7337__I0 _3640_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8370__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6465_ _3065_ _3069_ _3071_ _3072_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__5899__I0 mod.Data_Mem.F_M.MRAM\[4\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8204_ _0305_ net1 mod.Data_Mem.F_M.MRAM\[12\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_106_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7938__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5416_ _2065_ _2075_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_134_759 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5512__A2 mod.Data_Mem.F_M.MRAM\[30\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6396_ _2092_ _3005_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_161_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8135_ mod.Data_Mem.F_M.out_data\[45\] net2 net1 mod.Arithmetic.CN.I_in\[45\] vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_5347_ mod.Data_Mem.F_M.MRAM\[791\]\[6\] mod.Data_Mem.F_M.MRAM\[788\]\[6\] mod.Data_Mem.F_M.MRAM\[789\]\[6\]
+ mod.Data_Mem.F_M.MRAM\[790\]\[6\] _1829_ _2009_ _2010_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_82_1046 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8066_ _0275_ net1 mod.Data_Mem.F_M.MRAM\[21\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_102_645 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5278_ _1514_ _1942_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__4079__A2 _0708_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_102_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7017_ _3239_ _3450_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_75_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4229_ _0839_ _0904_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_75_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5399__I _2059_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6225__B1 mod.Data_Mem.F_M.MRAM\[15\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7919_ _0145_ net1 mod.Data_Mem.F_M.MRAM\[0\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_24_640 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_145_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_1153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_278 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6528__A1 _2626_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_51_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7576__I0 _3749_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_169_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_169_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7119__I _3252_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6023__I _2388_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_165_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_152_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5503__A2 _2142_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_93_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_98_1020 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_1015 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4490__A2 _1082_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_713 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8243__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5102__I _1701_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_1086 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2050 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2061 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2072 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2083 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4242__A2 mod.Arithmetic.ACTI.x\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_1204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8560__D _0064_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2094 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1360 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6519__A1 _3120_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1371 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7567__I0 _3731_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1382 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5990__A2 _2609_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_159_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1393 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_148_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__8393__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4580_ _1251_ _1250_ _1136_ _1017_ _1252_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_155_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_726 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6250_ _2212_ _1627_ _2864_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_115_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5201_ _1757_ mod.Data_Mem.F_M.MRAM\[15\]\[3\] mod.Data_Mem.F_M.MRAM\[31\]\[3\] _1721_
+ _1866_ _1867_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_42_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4388__I _0632_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6181_ _2687_ _2795_ _2796_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5132_ _1669_ _1799_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_96_120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5258__A1 _1704_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6309__S _2723_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5063_ _1602_ _1730_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_97_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5213__S _1877_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4014_ mod.Arithmetic.CN.I_in\[20\] _0691_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_65_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_168_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5965_ _1627_ _2143_ _2145_ _2585_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_7704_ mod.Data_Mem.F_M.MRAM\[793\]\[4\] _3846_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4916_ _1584_ _1585_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_5896_ _2510_ _2514_ _2516_ _2517_ _2518_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_33_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5981__A2 _2598_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7635_ _3811_ _0505_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4847_ mod.Data_Mem.F_M.MRAM\[19\]\[0\] mod.Data_Mem.F_M.MRAM\[18\]\[0\] _1515_ _1516_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_147_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7566_ _3769_ _0478_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4778_ _1309_ _1317_ _1448_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_88_1200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_107_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6517_ _3049_ _2329_ _3050_ _2578_ _2580_ _2496_ _3121_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_106_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5682__I _2069_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7497_ _3725_ mod.Data_Mem.F_M.MRAM\[781\]\[4\] _3726_ _3727_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_49_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_106_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_1119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6448_ _3004_ _3054_ _3055_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5497__A1 _1686_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8116__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_164_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_106_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6379_ _2886_ _2985_ _2988_ _2989_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_88_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7603__S _3787_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8118_ mod.Data_Mem.F_M.out_data\[28\] net2 net1 mod.Arithmetic.CN.I_in\[28\] vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_130_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_569 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_88_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_87_153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_987 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_8049_ _0258_ net1 mod.Data_Mem.F_M.MRAM\[1\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_75_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8266__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4847__I1 mod.Data_Mem.F_M.MRAM\[18\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_1152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_584 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_71_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7797__I0 _3319_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_31_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_169_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_169_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_1013 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_169_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6221__I0 mod.Data_Mem.F_M.MRAM\[1\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_32_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5724__A2 _2156_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5592__I _1811_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_153_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_125_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5488__B2 _2133_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_106_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_1030 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_610 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7513__S _3734_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_429 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_117_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_773 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7312__I _3622_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5335__S1 _1882_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_152_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5660__A1 _2290_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7788__I0 _3306_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_90_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4215__A2 _0834_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5750_ _1595_ _1500_ _2375_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_76_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1190 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4701_ _1370_ _1247_ _1371_ _1372_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_5681_ _2305_ _2310_ _0051_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_31_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_7420_ _3683_ _0418_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4632_ mod.Arithmetic.CN.I_in\[37\] _1214_ _1303_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_129_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5715__A2 _2337_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_159_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8139__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4563_ _1111_ _1120_ _1233_ _1235_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_7351_ mod.Data_Mem.F_M.MRAM\[772\]\[0\] _3649_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_128_394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6302_ _2866_ _2914_ _0068_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_7282_ _3297_ _3604_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_4494_ _1052_ _1074_ _1166_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6233_ _1802_ _1832_ _2846_ _2847_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_131_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6140__A2 _2755_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8289__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5007__I _1514_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4151__A1 _0652_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_930 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_83_1163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6164_ _1555_ _1702_ _1703_ _1566_ _2780_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_462 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4846__I _1514_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5115_ _1518_ _1782_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_974 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_924 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_985 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_84_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6095_ _2196_ _1604_ _2712_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5046_ _1578_ _1714_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_85_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2808 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_713 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2819 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_66_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_168_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6997_ _3437_ _0241_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_25_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5948_ _1778_ mod.Data_Mem.F_M.MRAM\[3\]\[4\] _2569_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__5954__A2 _1870_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_40_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5879_ mod.Data_Mem.F_M.MRAM\[788\]\[3\] mod.Data_Mem.F_M.MRAM\[789\]\[3\] _2161_
+ _2501_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_7618_ _3749_ mod.Data_Mem.F_M.MRAM\[787\]\[2\] _3801_ _3802_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_166_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5706__A2 _2329_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7549_ _3232_ _3298_ _3758_ _3759_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_4_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_162_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4142__A1 _0812_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_322 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_816 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_773 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_102_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6176__C _2374_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5642__A1 _2264_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_178 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_1001 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_1045 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5945__A2 _2137_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_251 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_284 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_158_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_33_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_9_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_832 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8431__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_1125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6367__B _2873_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4684__A2 _1354_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8581__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_819 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4436__A2 _0995_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6881__I mod.Data_Mem.F_M.MRAM\[4\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_1210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6920_ _3227_ _3386_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_165_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6851_ mod.Data_Mem.F_M.MRAM\[779\]\[1\] _3348_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6189__A2 mod.Data_Mem.F_M.MRAM\[6\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5802_ _2425_ mod.Data_Mem.F_M.MRAM\[785\]\[1\] _2426_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_50_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3994_ _0649_ _0670_ _0671_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__5936__A2 _2556_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6782_ _3302_ _3303_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_8521_ _0025_ net1 mod.Data_Mem.F_M.out_data\[49\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5733_ _1681_ _2358_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_8452_ _0548_ net1 mod.Data_Mem.F_M.MRAM\[794\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_148_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5664_ _1686_ _2295_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_7403_ mod.Data_Mem.F_M.MRAM\[775\]\[2\] _3675_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4615_ _1205_ _1218_ _1286_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_8383_ _0479_ net1 mod.Data_Mem.F_M.MRAM\[784\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5595_ mod.Data_Mem.F_M.MRAM\[29\]\[4\] _2226_ _2227_ mod.Data_Mem.F_M.MRAM\[28\]\[4\]
+ _2231_ _2232_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XFILLER_135_128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_832 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7217__I _3561_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_11_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_4546_ _1207_ _1212_ _1217_ _1218_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
X_7334_ _3638_ mod.Data_Mem.F_M.MRAM\[771\]\[1\] _3636_ _3639_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_144_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_504 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_898 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7265_ mod.Data_Mem.F_M.MRAM\[5\]\[0\] _3595_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6113__A2 mod.Data_Mem.F_M.MRAM\[3\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4477_ _0725_ _0716_ _0816_ _0972_ _1149_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_2
XFILLER_104_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7161__I1 mod.Data_Mem.F_M.MRAM\[12\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6216_ _2797_ _2803_ _2830_ _2374_ _0066_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_7196_ _3308_ _3555_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_98_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_1050 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5872__A1 _2085_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_782 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6147_ _2713_ _2763_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_100_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_38_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_771 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_782 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_793 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6078_ _2684_ _2688_ _1726_ _2694_ _2695_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_57_167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5624__A1 _2256_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5029_ _1674_ _1696_ _1558_ _1697_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_2605 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2616 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2627 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2638 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2649 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1904 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1915 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8304__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1926 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1937 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1948 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_13_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_81_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1959 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5200__I _1669_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_1130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_1073 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8454__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_167_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5356__B _1775_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7127__I _3512_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5155__A3 _1820_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_5_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5560__B1 _2195_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_163_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_898 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_79_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_846 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4115__A1 mod.Arithmetic.ACTI.x\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4115__B2 mod.Arithmetic.ACTI.x\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_50 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_27_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_1180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6187__B _1965_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_150_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_95_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xtiny_user_project_101 la_data_out[22] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_112 la_data_out[33] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_123 la_data_out[44] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_134 la_data_out[55] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XANTENNA__6407__A3 _3015_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xtiny_user_project_145 user_irq[2] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_48_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_1107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xtiny_user_project_156 wbs_dat_o[9] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_36_307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8097__RN net2 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5615__A1 _2225_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4418__A2 _1090_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5615__B2 _2177_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xtiny_user_project_167 wbs_dat_o[20] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_91_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xtiny_user_project_178 wbs_dat_o[31] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_64_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5091__A2 mod.Data_Mem.F_M.MRAM\[31\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5218__I1 _1876_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6966__I1 mod.Data_Mem.F_M.MRAM\[15\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6040__A1 _2549_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_32_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_1162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7238__S _3579_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_157_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6343__A2 _2952_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4400_ _1067_ _1072_ _1073_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5380_ mod.Data_Mem.F_M.MRAM\[773\]\[7\] mod.Data_Mem.F_M.MRAM\[772\]\[7\] _1906_
+ _2042_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_154_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_126_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4331_ _0911_ _0919_ _1005_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_114_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7143__I1 mod.Data_Mem.F_M.MRAM\[19\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7050_ _3456_ mod.Data_Mem.F_M.MRAM\[1\]\[4\] _3469_ _3472_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__4106__B2 _0781_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4262_ _0865_ _0936_ _0937_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__7971__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_80_1111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6001_ _1681_ _2620_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_68_911 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5854__A1 _2475_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4657__A2 _1212_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_933 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4193_ _0639_ _0811_ _0868_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_132_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_966 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_977 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8327__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8088__RN net2 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_1199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5606__A1 _1940_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7952_ _0178_ net1 mod.Data_Mem.F_M.MRAM\[769\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_55_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_1040 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6903_ _3228_ mod.Data_Mem.F_M.MRAM\[13\]\[0\] _3376_ _3377_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_7883_ _0109_ net1 mod.Data_Mem.F_M.MRAM\[26\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__5209__I1 mod.Data_Mem.F_M.MRAM\[4\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6834_ _3240_ mod.Data_Mem.F_M.MRAM\[769\]\[1\] _3337_ _3339_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__8477__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6031__A1 _2506_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6765_ _3289_ _0157_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_23_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6582__A2 _3179_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3977_ _0653_ _0654_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__7148__S _3525_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4999__C _1616_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8504_ _0008_ net1 mod.Data_Mem.F_M.out_data\[64\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__4593__A1 _0786_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5716_ _2342_ _0054_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__5790__B1 _2412_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_149_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6696_ _3246_ mod.Data_Mem.F_M.MRAM\[28\]\[3\] _3237_ _3247_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__6709__I1 mod.Data_Mem.F_M.MRAM\[28\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8435_ _0531_ net1 mod.Data_Mem.F_M.MRAM\[792\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__6987__S _3428_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_163_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5647_ _2168_ _2278_ _2279_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__4345__A1 _0617_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8366_ _0462_ net1 mod.Data_Mem.F_M.MRAM\[782\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5578_ _1493_ _2216_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_3_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_1082 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7317_ _1765_ _3626_ _3628_ _0370_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__6786__I _3305_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5690__I _2096_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4529_ _1198_ _1199_ _1200_ _1201_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__7134__I1 mod.Data_Mem.F_M.MRAM\[19\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8297_ _0393_ net1 mod.Data_Mem.F_M.MRAM\[773\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_46_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_868 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7248_ mod.Data_Mem.F_M.MRAM\[31\]\[0\] _3293_ _3585_ _3586_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_132_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_59_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5845__A1 _2425_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7179_ mod.Data_Mem.F_M.MRAM\[22\]\[4\] _3545_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_86_730 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_432 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3103 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8079__RN net2 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3114 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_796 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3125 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3136 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3147 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2402 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2413 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3158 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5073__A2 _1739_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3169 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2424 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2435 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_73_468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2446 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1701 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2457 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1712 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2468 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1723 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_57_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2479 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_157_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_41_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_1157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1745 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_546 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1756 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1048 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6022__A1 _2587_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1767 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1778 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1789 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_139_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_108_640 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4336__A1 _0642_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7994__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_108_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4887__A2 _1555_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_155_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5306__S _1515_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_1117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_816 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_111_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4639__A2 mod.Arithmetic.CN.I_in\[22\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xtiny_user_project_40 io_oeb[29] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_51 io_out[2] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_77_752 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xtiny_user_project_62 io_out[13] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_49_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xtiny_user_project_73 io_out[32] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_65_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtiny_user_project_84 la_data_out[5] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_92_711 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_796 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtiny_user_project_95 la_data_out[16] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_37_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6261__A1 _2872_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_80_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_162_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2980 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_32_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4880_ _1504_ _1549_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_72_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2991 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6939__I1 mod.Data_Mem.F_M.MRAM\[14\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6013__A1 _2549_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6564__A2 _2655_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6550_ _2728_ mod.Data_Mem.F_M.MRAM\[1\]\[7\] _3152_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_125_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5501_ _2144_ mod.Data_Mem.F_M.MRAM\[31\]\[5\] _2145_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_72_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_145_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6316__A2 _1957_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6481_ _2264_ mod.Data_Mem.F_M.MRAM\[781\]\[3\] _3087_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_8220_ _0321_ net1 mod.Data_Mem.F_M.MRAM\[29\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__4327__A1 _0993_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_161_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5432_ _2086_ _2087_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5524__B1 _2160_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4878__A2 _1532_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5363_ _1835_ _2025_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_8151_ mod.Data_Mem.F_M.out_data\[61\] net2 net1 mod.Arithmetic.CN.I_in\[61\] vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_99_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7102_ mod.Data_Mem.F_M.MRAM\[23\]\[6\] _3498_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_99_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4314_ _0979_ _0987_ _0988_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_99_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8082_ _0282_ net1 mod.Data_Mem.F_M.MRAM\[23\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5294_ mod.Data_Mem.F_M.MRAM\[771\]\[5\] mod.Data_Mem.F_M.MRAM\[770\]\[5\] _1783_
+ _1958_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_114_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7033_ _3460_ mod.Data_Mem.F_M.MRAM\[18\]\[6\] _3457_ _3461_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4245_ _0911_ _0914_ _0919_ _0920_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_45_1061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_730 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_28_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4176_ _0819_ _0851_ _0852_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_67_251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5055__A2 _1699_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6252__A1 _2534_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_167_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_55_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_788 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7935_ _0161_ net1 mod.Data_Mem.F_M.MRAM\[799\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__7867__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1019 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4802__A2 _1457_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7866_ _0092_ net1 mod.Data_Mem.F_M.MRAM\[11\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_35_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6004__A1 _2588_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6817_ _3327_ _0171_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4015__B1 _0680_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7797_ _3319_ mod.Data_Mem.F_M.MRAM\[798\]\[6\] _3894_ _3897_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_51_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6555__A2 _3153_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_1021 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4566__A1 _0618_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6748_ _3253_ mod.Data_Mem.F_M.MRAM\[0\]\[5\] _3279_ _3281_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_50_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5618__C _2251_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6679_ mod.DMen_reg2 _3233_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_104_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5515__B1 _2156_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8418_ _0514_ net1 mod.Data_Mem.F_M.MRAM\[790\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__4318__B2 _0933_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_164_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_151_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_8349_ _0445_ net1 mod.Data_Mem.F_M.MRAM\[780\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__7405__I mod.Data_Mem.F_M.MRAM\[775\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5818__A1 _2283_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_23 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_63_1161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6491__A1 _2728_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_914 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_785 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_755 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2210 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2221 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2232 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2243 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2254 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2265 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1520 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2276 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1531 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2287 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1542 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_60 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_14_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1553 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7043__I0 _3450_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2298 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_71 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_41_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_82 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1575 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__6546__A2 _2341_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1586 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1597 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4557__A1 mod.Arithmetic.CN.I_in\[53\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8022__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_168_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_10_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_571 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__4309__A1 _0650_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_6_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8172__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4939__I _1607_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5263__C _1629_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_155_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_116_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4875__S _1543_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4030_ mod.Arithmetic.CN.I_in\[10\] _0707_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__6482__A1 _2475_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_755 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6234__A1 _2723_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5981_ _2596_ _2598_ _2600_ _2397_ _2601_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_18_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5588__A3 _2093_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7720_ mod.Data_Mem.F_M.MRAM\[794\]\[4\] _3854_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_52_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_1021 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_1190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4932_ _1600_ _1601_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_45_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_162_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7651_ _3819_ _0513_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4863_ mod.Data_Mem.F_M.MRAM\[22\]\[0\] _1511_ _1516_ _1520_ _1527_ _1531_ _1532_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_33_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6537__A2 _2210_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6602_ _3191_ _0092_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_21_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4548__A1 _1122_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7582_ _3778_ mod.Data_Mem.F_M.MRAM\[785\]\[4\] _3779_ _3780_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_32_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4794_ _1423_ _1331_ _1464_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_6533_ _2522_ mod.Data_Mem.F_M.MRAM\[0\]\[6\] _2102_ _3136_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__8515__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_158_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6464_ _2831_ _3070_ _2073_ _3071_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_133_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8203_ _0304_ net1 mod.Data_Mem.F_M.MRAM\[12\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__5899__I1 mod.Data_Mem.F_M.MRAM\[5\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4849__I _1517_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5415_ _2073_ _2074_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_86_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6395_ _2698_ _3004_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_82_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8134_ mod.Data_Mem.F_M.out_data\[44\] net2 net1 mod.Arithmetic.CN.I_in\[44\] vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_88_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5346_ _2008_ _2009_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_88_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_114_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8065_ _0274_ net1 mod.Data_Mem.F_M.MRAM\[21\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5277_ _1940_ _1941_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__7161__S _3534_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6473__A1 _3014_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7016_ _3449_ _0248_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4228_ _0901_ _0902_ _0903_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_101_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_68_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_56_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4159_ _0830_ _0834_ _0835_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_46_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6225__A1 _2217_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6225__B2 _2319_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_788 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7918_ _0144_ net1 mod.Data_Mem.F_M.MRAM\[0\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__8045__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4787__A1 _0624_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_168_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_1116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_1165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7849_ mod.Data_Mem.F_M.MRAM\[9\]\[3\] _3927_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6528__A2 _3129_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_169_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_62_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4539__A1 _1209_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_11_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8195__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5339__I0 mod.Data_Mem.F_M.MRAM\[769\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_65_1201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_1212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_79_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_911 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_133_771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6839__I0 _3246_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6464__A1 _2831_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_498 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_427 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5814__I1 mod.Data_Mem.F_M.MRAM\[783\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2040 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2051 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2062 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2073 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2084 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1350 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2095 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1361 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_1216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1372 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8538__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7567__I1 mod.Data_Mem.F_M.MRAM\[784\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1394 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_35_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_1009 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7045__I _3465_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5200_ _1669_ _1866_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4702__A1 _0643_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6180_ mod.Data_Mem.F_M.MRAM\[781\]\[2\] _2200_ _2202_ mod.Data_Mem.F_M.MRAM\[780\]\[2\]
+ _2794_ _2795_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_69_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5131_ _1759_ _1796_ _1797_ _1558_ _1798_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_97_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5258__A2 _1922_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5062_ _1537_ _1729_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_96_154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_677 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_1020 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_85_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4013_ mod.Arithmetic.I_out\[76\] _0690_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_38_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_65_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8068__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6207__A1 _2708_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_1116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_53_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4769__A1 _0624_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5964_ _2558_ _2580_ _2583_ _2584_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__7007__I0 _3403_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7703_ _3845_ _0539_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4915_ _1564_ _1584_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_61_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5895_ _2116_ _2517_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_33_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_166_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_7634_ mod.Data_Mem.F_M.MRAM\[788\]\[1\] _3811_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4846_ _1514_ _1515_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__7905__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5194__A1 _1721_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7565_ _3729_ mod.Data_Mem.F_M.MRAM\[784\]\[6\] _3759_ _3769_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_165_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4777_ _1297_ _1445_ _1446_ _1447_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_88_1212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6516_ _3115_ _3116_ _3119_ _2434_ _3120_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_162_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7496_ _3719_ _3726_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_107_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4579__I _1061_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6447_ _3005_ _2292_ _3006_ _2466_ _2469_ _3023_ _3054_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XANTENNA__5497__A2 mod.Data_Mem.F_M.MRAM\[799\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_161_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6378_ _2733_ _2986_ _2987_ _2988_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_103_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8117_ mod.Data_Mem.F_M.out_data\[27\] net2 net1 mod.Arithmetic.CN.I_in\[27\] vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_88_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5912__B _2533_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_730 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5329_ _1872_ _1991_ _1863_ _1992_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_103_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_432 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8048_ _0257_ net1 mod.Data_Mem.F_M.MRAM\[1\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_88_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_1164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_1_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_84_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_95_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_714 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_894 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_43_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_106_1025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_975 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_157_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6382__B1 _2991_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5873__I _2101_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_152_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_125_535 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_156_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5314__S _1568_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8210__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6437__A1 _2312_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5660__A2 _2125_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_574 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_500 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8360__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8571__D _0075_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7928__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6372__C _2078_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_717 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1180 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4700_ _1242_ _1246_ _1371_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_148_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1191 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_1046 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_290 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5680_ _2306_ _2309_ _2310_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_30_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4631_ _1301_ _1302_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__5176__A1 _1840_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_147_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7350_ _3648_ _0383_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5971__I0 mod.Data_Mem.F_M.MRAM\[2\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4562_ _1111_ _1120_ _1233_ _1234_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_144_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6301_ _2868_ _2900_ _2913_ _2914_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_7281_ _3292_ _3603_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6125__B1 _2737_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4493_ _1049_ _1163_ _1164_ _1165_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_143_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_568 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5479__A2 _2124_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6232_ _2714_ _2846_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_83_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4151__A2 _0826_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6163_ _2707_ _2779_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_98_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_931 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_942 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5224__S _1588_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_1175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6428__A1 _1933_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_964 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7476__I0 _3615_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5114_ _1778_ mod.Data_Mem.F_M.MRAM\[791\]\[2\] _1780_ _1781_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_98_997 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_975 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6094_ _2326_ mod.Data_Mem.F_M.MRAM\[790\]\[0\] mod.Data_Mem.F_M.MRAM\[791\]\[0\]
+ _2116_ _2711_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_986 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_997 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5100__A1 _1707_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5045_ _1526_ _1713_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_38_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4454__A3 _0914_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2809 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_84_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4862__I _1530_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6055__S _1769_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6996_ _3393_ mod.Data_Mem.F_M.MRAM\[17\]\[1\] _3435_ _3437_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_80_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5947_ _2102_ _2568_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_90_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_167_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5878_ _2499_ _2500_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_90_1157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7617_ _3797_ _3801_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__6789__I net6 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5167__A1 _1764_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4829_ _1497_ _1498_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_21_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4914__A1 _1575_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7548_ _3420_ _3758_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_88_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7479_ _3715_ _0445_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_88_1075 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8233__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8510__188 net188 vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_134_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_89_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_538 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_942 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_1204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3941__I _0618_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_430 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6419__A1 _2626_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8383__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_5_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_500 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_241 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_252 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_285 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__5158__A1 _1805_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_158_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7524__S _3739_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_739 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_165_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_398 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5330__A1 mod.Data_Mem.F_M.MRAM\[31\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_67_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_94_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_820 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5778__I _2402_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6850_ _3347_ _0184_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_39_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5801_ _1636_ _2425_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__8106__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6781_ net4 _3302_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_50_536 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3993_ _0652_ _0657_ _0669_ _0670_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
X_8520_ _0024_ net1 mod.Data_Mem.F_M.out_data\[48\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5732_ _2356_ _2357_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_50_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_8451_ _0547_ net1 mod.Data_Mem.F_M.MRAM\[794\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_31_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5663_ _2135_ mod.Data_Mem.F_M.MRAM\[29\]\[2\] _2294_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__8256__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7402_ _3674_ _0409_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4614_ _1283_ _1195_ _1284_ _1285_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_8382_ _0478_ net1 mod.Data_Mem.F_M.MRAM\[784\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__4747__I1 mod.Arithmetic.CN.I_in\[70\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5594_ _2228_ _2230_ _2231_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_116_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7333_ _3302_ _3638_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4372__A2 _1024_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4545_ _1213_ _1216_ _1217_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__5018__I _1594_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_7264_ _3594_ _0351_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4476_ _1031_ _1032_ _1034_ _1148_ mod.P3.Res\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_131_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4857__I _1525_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6215_ _1800_ _2818_ _2823_ _2829_ _2743_ _2830_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XANTENNA__5321__A1 _1966_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7195_ _3554_ _0322_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_131_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6146_ _2761_ _1637_ _2762_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_1062 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_761 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6077_ _2087_ _2690_ _2693_ _2694_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__5624__A2 mod.Data_Mem.F_M.MRAM\[797\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5028_ _1680_ _1684_ _1689_ _1694_ _1695_ _1651_ _1696_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XTAP_2606 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2617 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2628 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2639 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_166_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_26_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1905 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1916 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1927 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_717 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_54_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_41_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5388__A1 _1875_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1938 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1949 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6979_ _3426_ _0234_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_80_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7609__S _3786_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_1030 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3936__I _0613_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_166_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5935__I0 mod.Data_Mem.F_M.MRAM\[18\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_107_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_135_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_162_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6468__B _3031_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_398 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5312__A1 _1622_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6360__I0 _2246_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_1001 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_603 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_1023 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_1192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_89_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xtiny_user_project_102 la_data_out[23] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_62_1056 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6982__I _3422_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xtiny_user_project_113 la_data_out[34] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_48_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xtiny_user_project_124 la_data_out[45] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XANTENNA__6499__S0 _2270_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xtiny_user_project_135 la_data_out[56] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_146 wbs_ack_o vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_76_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5615__A2 _2246_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_617 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_1119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xtiny_user_project_157 wbs_dat_o[10] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_168 wbs_dat_o[21] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_48_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8129__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_149_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_91_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_801 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5218__I2 _1878_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8279__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4007__I mod.Arithmetic.CN.I_in\[17\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_1174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_160_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5551__A1 _2186_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7254__S _3585_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4330_ _0921_ _0926_ _1003_ _1004_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_4_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_1035 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_113_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_158_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5303__A1 mod.Data_Mem.F_M.MRAM\[15\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6351__I0 _1994_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4261_ _0866_ _0886_ _0935_ _0936_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_87_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_901 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6000_ _1778_ _2619_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_140_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4192_ _0623_ _0656_ _0820_ _0835_ _0867_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
XANTENNA_input2_I io_in[9] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_94_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_606 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7951_ _0177_ net1 mod.Data_Mem.F_M.MRAM\[769\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_94_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_285 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6902_ _3375_ _3376_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_82_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7882_ _0108_ net1 mod.Data_Mem.F_M.MRAM\[26\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_51_801 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_36_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7603__I0 _3778_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6833_ _3338_ _0176_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_50_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6031__A2 mod.Data_Mem.F_M.MRAM\[788\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6764_ mod.Data_Mem.F_M.MRAM\[8\]\[5\] _3289_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_11_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3976_ _0616_ _0653_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_8503_ _0007_ net1 mod.Data_Mem.F_M.out_data\[79\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5715_ _2082_ _2337_ _2341_ _2306_ _2342_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__5790__A1 _1491_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6695_ _3245_ _3246_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_148_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5790__B2 _2414_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8434_ _0530_ net1 mod.Data_Mem.F_M.MRAM\[792\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5646_ _2274_ _2276_ _2277_ _2278_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_164_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_8365_ _0461_ net1 mod.Data_Mem.F_M.MRAM\[782\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__5542__A1 _2180_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4345__A2 _1017_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5577_ _2214_ mod.Data_Mem.F_M.MRAM\[31\]\[3\] _2215_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_105_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_1181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_163_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7316_ _3612_ _3623_ _3628_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_144_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4528_ _1108_ _1140_ _1200_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_102_1094 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8296_ _0392_ net1 mod.Data_Mem.F_M.MRAM\[773\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_46_1007 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_160_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7295__A1 _3555_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7247_ _3584_ _3585_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__6342__I0 _2015_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4459_ _1125_ _1131_ _1132_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_120_806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_104_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_7178_ _3544_ _0315_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_58_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6129_ _2619_ mod.Data_Mem.F_M.MRAM\[783\]\[1\] mod.Data_Mem.F_M.MRAM\[782\]\[1\]
+ _2089_ _2745_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3104 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_926 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3115 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3126 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3137 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3148 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2403 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3159 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2414 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2425 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2436 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4281__A1 _0877_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1702 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2447 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8421__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2458 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1713 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2469 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1724 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1735 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6558__B1 _2663_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1746 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6022__A2 mod.Data_Mem.F_M.MRAM\[5\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1757 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7339__S _3636_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1768 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_878 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1779 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8571__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_167_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4336__A2 mod.Arithmetic.ACTI.x\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5533__A1 mod.Data_Mem.F_M.MRAM\[797\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5881__I _2376_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_163_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_155_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6089__A2 _1542_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_150_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_123_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4639__A3 _0678_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_462 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtiny_user_project_30 io_oeb[19] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_41 io_oeb[30] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_52 io_out[3] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_39_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xtiny_user_project_63 io_out[14] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_7_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_77_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xtiny_user_project_74 io_out[33] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_85 la_data_out[6] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_77_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xtiny_user_project_96 la_data_out[17] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_36_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__6261__A2 _1876_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6217__I _2107_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_789 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2970 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2981 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2992 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_355 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4024__A1 _0696_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5072__I0 mod.Data_Mem.F_M.MRAM\[3\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5500_ _2059_ _2144_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_9_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6480_ _3031_ _3085_ _3047_ _3086_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_146_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6887__I mod.Data_Mem.F_M.MRAM\[4\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5431_ _1549_ _2086_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_65_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4327__A2 _0999_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5524__A1 mod.Data_Mem.F_M.MRAM\[29\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5524__B2 _2164_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_145_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_983 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_126_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8150_ mod.Data_Mem.F_M.out_data\[60\] net2 net1 mod.Arithmetic.CN.I_in\[60\] vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_5362_ mod.Data_Mem.F_M.MRAM\[1\]\[7\] mod.Data_Mem.F_M.MRAM\[0\]\[7\] _1879_ _2024_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_99_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7101_ _3497_ _0285_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_142_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4313_ _0982_ _0986_ _0987_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_8081_ _0281_ net1 mod.Data_Mem.F_M.MRAM\[23\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_82_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5293_ _1954_ _1955_ _1956_ _1957_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_99_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7032_ _3255_ _3460_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_113_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4244_ _0916_ _0918_ _0919_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__5383__S0 _2044_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_1021 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_101_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4175_ _0823_ _0850_ _0851_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__8444__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_572 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7934_ _0160_ net1 mod.Data_Mem.F_M.MRAM\[799\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1009 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_70_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7865_ _0091_ net1 mod.Data_Mem.F_M.MRAM\[11\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__8594__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_169_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4870__I _1538_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6816_ mod.Data_Mem.F_M.MRAM\[789\]\[3\] _3327_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_24_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_7796_ _3896_ _0581_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_17_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6998__S _3435_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6747_ _3280_ _0148_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4566__A2 mod.Arithmetic.CN.I_in\[68\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3959_ _0635_ _0636_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_149_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7992__RN net2 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6678_ _3231_ _3232_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__5515__A1 _2119_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5629_ _2094_ _2261_ _2262_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_8417_ _0513_ net1 mod.Data_Mem.F_M.MRAM\[790\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_118_950 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5515__B2 _2133_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8348_ _0444_ net1 mod.Data_Mem.F_M.MRAM\[780\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_145_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_964 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_105_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8279_ _0375_ net1 mod.Data_Mem.F_M.MRAM\[770\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_132_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5818__A2 mod.Data_Mem.F_M.MRAM\[773\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5374__S0 _1844_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_59_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_120_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6491__A2 mod.Data_Mem.F_M.MRAM\[1\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5142__S _1510_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2200 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4981__S _1509_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2211 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2222 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2233 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2244 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2255 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1510 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2266 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2277 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1532 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2288 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_50 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1543 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_951 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7043__I1 mod.Data_Mem.F_M.MRAM\[1\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2299 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_61 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_14_344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1554 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_72 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1565 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_83 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_70_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7961__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_94 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1587 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_42_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_1111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1598 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4557__A2 _1114_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7983__RN net2 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_70_1188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5506__A1 _1677_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4309__A2 mod.Arithmetic.CN.I_in\[43\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8317__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5317__S _1568_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_1040 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_430 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5116__I _1567_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8467__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_151_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_96_325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_859 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8574__D _0078_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_1213 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8160__RN net2 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_926 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_37_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_65_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6234__A2 _1830_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5980_ _2343_ mod.Data_Mem.F_M.MRAM\[772\]\[5\] _2599_ _2600_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_24_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_64_288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4931_ _1523_ _1600_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5993__A1 _2588_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7650_ mod.Data_Mem.F_M.MRAM\[790\]\[1\] _3819_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4862_ _1530_ _1531_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_36_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_675 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6537__A3 _2636_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6601_ mod.Data_Mem.F_M.MRAM\[11\]\[4\] _3191_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_20_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5745__A1 _2366_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7581_ _3772_ _3779_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_4793_ _1422_ _1462_ _1463_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6532_ _2061_ mod.Data_Mem.F_M.MRAM\[1\]\[6\] _3135_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_6463_ _3005_ _2298_ _3009_ _2487_ _2491_ _3023_ _3070_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_118_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8202_ _0087_ net2 net1 mod.I_addr\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_5414_ _1725_ _2073_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_134_739 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5899__I2 mod.Data_Mem.F_M.MRAM\[20\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6170__A1 _2196_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6394_ _1724_ _3003_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_86_1140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_249 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_8133_ mod.Data_Mem.F_M.out_data\[43\] net2 net1 mod.Arithmetic.CN.I_in\[43\] vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_86_1162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5345_ _1914_ _2008_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_86_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_975 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_1184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8064_ _0273_ net1 mod.Data_Mem.F_M.MRAM\[21\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_102_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5276_ _1573_ _1940_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_7015_ _3445_ mod.Data_Mem.F_M.MRAM\[18\]\[0\] _3448_ _3449_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__4865__I mod.Data_Mem.F_M.src\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4227_ _0890_ _0900_ _0902_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_102_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8151__RN net2 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4158_ _0832_ _0833_ _0834_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_110_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4086__B _0710_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6225__A2 mod.Data_Mem.F_M.MRAM\[14\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4089_ _0746_ _0766_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_83_575 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7984__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_1100 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7917_ _0143_ net1 mod.Data_Mem.F_M.MRAM\[10\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_70_225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4787__A2 _1456_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5984__A1 _2424_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_951 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_145_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_169_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7848_ _3926_ _0602_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_23_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_1128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7779_ _3886_ _0574_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_168_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_125_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5339__I1 mod.Data_Mem.F_M.MRAM\[768\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3944__I _0621_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_164_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6161__A1 _2681_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_513 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_975 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_133_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6839__I1 mod.Data_Mem.F_M.MRAM\[769\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5347__S0 _1829_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8142__RN net2 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6464__A2 _3070_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__4475__A1 _1031_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_19_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2030 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2041 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5975__A1 _2531_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2052 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_61_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2063 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2074 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1340 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2085 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2096 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1362 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1373 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1384 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1395 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_156_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_157_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4702__A2 mod.Arithmetic.CN.I_in\[70\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_761 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5130_ mod.Data_Mem.F_M.MRAM\[799\]\[2\] _1775_ _1797_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_123_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_28_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__8133__RN net2 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5061_ _1728_ _0001_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_4012_ _0680_ _0681_ _0682_ _0683_ _0686_ _0688_ _0689_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai222_4
XFILLER_84_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_168_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_52_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5963_ _2397_ _2581_ _2582_ _2583_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__5966__A1 _2579_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4769__A2 _1134_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7007__I1 mod.Data_Mem.F_M.MRAM\[17\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7702_ mod.Data_Mem.F_M.MRAM\[793\]\[3\] _3845_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6405__I _2100_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4914_ _1575_ _1582_ _1583_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_33_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_80_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5894_ _2511_ _1846_ _2515_ _2516_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_7633_ _3810_ _0504_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5718__A1 _2343_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4845_ _1513_ _1514_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_60_291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7564_ _3768_ _0477_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4776_ _1300_ _1321_ _1446_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6515_ _3060_ _2591_ _2592_ _3020_ _3118_ _3119_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
X_7495_ _3311_ _3725_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_101_1126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_119_588 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_146_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_739 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_6446_ _3053_ _0073_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__7191__I0 _3527_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_162_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6377_ _2872_ _2043_ _2987_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_121_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_8116_ mod.Data_Mem.F_M.out_data\[26\] net2 net1 mod.Arithmetic.CN.I_in\[26\] vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_0_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5328_ _1987_ _1988_ _1989_ _1990_ _1881_ _1882_ _1991_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_102_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_87_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8047_ _0256_ net1 mod.Data_Mem.F_M.MRAM\[1\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_76_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8124__RN net2 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5259_ _1834_ _1921_ _1923_ _1642_ _1924_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__8012__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_169_1009 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_28_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_575 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4209__A1 mod.Arithmetic.CN.I_in\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8162__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5957__A1 _2534_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5957__B2 _2414_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3939__I _0616_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_169_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5709__A1 _2315_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_145_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7347__S _3643_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_156_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_132_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__6221__I2 mod.Data_Mem.F_M.MRAM\[3\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_987 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5375__B _1621_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4696__A1 _1134_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_133_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_753 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__8115__RN net2 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6437__A2 _2459_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8505__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_748 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_759 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5948__A1 _1778_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6996__I0 _3393_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4620__A1 _0828_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_163_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_1183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6748__I0 _3253_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1181 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1192 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7257__S _3590_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4630_ _1169_ _1183_ _1301_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__6373__A1 _1655_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5176__A2 mod.Data_Mem.F_M.MRAM\[775\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4561_ _1224_ _1232_ _1233_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_162_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_129_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_128_363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5971__I1 mod.Data_Mem.F_M.MRAM\[3\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6300_ _2703_ _2912_ _2913_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_7280_ _3602_ _0359_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6125__A1 _2696_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4492_ _1075_ _1076_ _1164_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__6125__B2 _2741_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6895__I mod.Data_Mem.F_M.MRAM\[4\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6231_ _2169_ _1837_ _2845_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_144_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_131_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8035__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6162_ _2769_ _2777_ _2778_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_910 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_943 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_69_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5113_ _1779_ mod.Data_Mem.F_M.MRAM\[790\]\[2\] _1780_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XTAP_954 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8106__RN net2 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_1187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_604 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_965 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6093_ _2705_ _2708_ _2709_ _2710_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XTAP_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_69_166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5304__I _1509_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_615 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4439__A1 _0650_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_987 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_998 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5044_ _1706_ _1711_ _1712_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_38_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8185__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5240__S _1836_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_501 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_168_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6563__C _2698_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_53_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6987__I0 _3403_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6995_ _3436_ _0240_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_25_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6135__I _1538_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_1201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5946_ _2283_ _2567_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_40_217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5877_ _2395_ _2499_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6739__I0 _3240_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_1169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4828_ _1493_ _1496_ _1497_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_7616_ _3800_ _0497_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6364__A1 _1585_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5167__A2 _1832_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7547_ _3757_ _0471_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4759_ _1418_ _1420_ _1428_ _1429_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XANTENNA__4914__A2 _1582_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_7478_ _3645_ mod.Data_Mem.F_M.MRAM\[780\]\[5\] _3713_ _3715_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_161_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_150_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6429_ _2620_ _1716_ _3036_ _3037_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_134_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8528__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6419__A2 _3027_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5214__I _1790_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_25_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6978__I0 _3395_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_16_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_898 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4602__A1 _0625_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_220 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_71_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__5884__I _2319_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_169_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_264 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_129_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_169_285 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_157_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_8_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_144_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__8058__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6107__A1 _2723_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_1116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5325__S _1873_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4669__A1 mod.Arithmetic.CN.I_in\[46\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5552__C _2191_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5330__A2 _1886_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5124__I _1790_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_572 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5618__B1 _1639_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_968 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4963__I _1628_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_47_394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_63_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5800_ _1612_ _2424_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_35_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6780_ _3301_ _0160_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_3992_ _0658_ _0668_ _0669_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_5731_ _2187_ _1499_ _2356_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_95_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5794__I _1517_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8450_ _0546_ net1 mod.Data_Mem.F_M.MRAM\[794\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_30_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6346__A1 _2876_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5662_ _2168_ _2292_ _2293_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4613_ _1165_ _1187_ _1284_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_7401_ mod.Data_Mem.F_M.MRAM\[775\]\[1\] _3674_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_8381_ _0477_ net1 mod.Data_Mem.F_M.MRAM\[784\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5593_ _1953_ mod.Data_Mem.F_M.MRAM\[31\]\[4\] mod.Data_Mem.F_M.MRAM\[30\]\[4\] _2229_
+ _2230_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_163_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4203__I _0877_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7332_ _3637_ _0376_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4544_ _1214_ _1215_ _1216_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_128_193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_1216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7263_ mod.Data_Mem.F_M.MRAM\[31\]\[7\] _3322_ _3590_ _3594_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4475_ _1031_ _1146_ _1147_ _1148_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_116_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6214_ _1898_ _2828_ _2829_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_116_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7194_ _3529_ mod.Data_Mem.F_M.MRAM\[29\]\[2\] _3553_ _3554_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_6145_ _1573_ _2761_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_751 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5609__B1 mod.Data_Mem.F_M.MRAM\[30\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_773 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_784 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6076_ mod.Data_Mem.F_M.MRAM\[781\]\[0\] _2692_ _2693_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_39_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_607 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4873__I _1541_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5027_ _1571_ _1695_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_39_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2607 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2618 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2629 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1906 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1917 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1928 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_504 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1939 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5388__A2 mod.Data_Mem.F_M.MRAM\[786\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_159_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6978_ _3395_ mod.Data_Mem.F_M.MRAM\[16\]\[2\] _3423_ _3426_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_1073 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_41_526 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_1020 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5929_ _2549_ mod.Data_Mem.F_M.MRAM\[772\]\[4\] _2550_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_167_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_146_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__8200__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6337__A1 _1635_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_155_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_8579_ _0595_ net1 mod.Instr_Mem.instruction\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__5935__I1 mod.Data_Mem.F_M.MRAM\[19\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7137__I0 _3456_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5560__A2 _2179_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_867 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8350__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7837__A1 _3913_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7918__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5312__A2 _1975_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6360__I1 _2249_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_1160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_773 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_615 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_76_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_946 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xtiny_user_project_103 la_data_out[24] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_103_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xtiny_user_project_114 la_data_out[35] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XANTENNA__6499__S1 _3083_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xtiny_user_project_125 la_data_out[46] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_76_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6484__B _3089_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xtiny_user_project_136 la_data_out[57] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_147 wbs_dat_o[0] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_158 wbs_dat_o[11] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_169 wbs_dat_o[22] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_64_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_29_383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_151_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_17_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_651 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5218__I3 _1880_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_846 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4051__A2 _0727_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6328__A1 _2752_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_73_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5926__I1 mod.Data_Mem.F_M.MRAM\[771\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_145_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7128__I0 _3445_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_92 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_125_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_113_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4260_ _0889_ _0903_ _0934_ _0935_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XANTENNA__6500__A1 _3083_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5303__A2 _1599_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6351__I1 _1995_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4191_ _0812_ _0817_ _0866_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_68_924 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7300__I0 _3569_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_1179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_55_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7950_ _0176_ net1 mod.Data_Mem.F_M.MRAM\[769\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_54_128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6901_ _3235_ _3371_ _3374_ _3375_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_78_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7881_ _0107_ net1 mod.Data_Mem.F_M.MRAM\[26\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_47_191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_169_1192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_982 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7603__I1 mod.Data_Mem.F_M.MRAM\[786\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6832_ _3228_ mod.Data_Mem.F_M.MRAM\[769\]\[0\] _3337_ _3338_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__8223__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6567__A1 _3003_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_165_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_62_194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6763_ _3288_ _0156_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_3975_ _0651_ mod.Arithmetic.CN.I_in\[32\] _0652_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_149_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_50_356 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8502_ _0006_ net1 mod.Data_Mem.F_M.out_data\[78\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5714_ _2316_ _2150_ _2338_ _2340_ _2341_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XANTENNA__6319__A1 _1603_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6694_ net6 _3245_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_31_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5790__A2 _2372_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8433_ _0529_ net1 mod.Data_Mem.F_M.MRAM\[792\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__8373__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5645_ _2270_ _2122_ _2277_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_108_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_8364_ _0460_ net1 mod.Data_Mem.F_M.MRAM\[782\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5576_ _2060_ _2214_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4868__I _1528_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4527_ _1108_ _1140_ _1199_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_7315_ _1709_ _3626_ _3627_ _0369_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_2_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_89_1193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8295_ _0391_ net1 mod.Data_Mem.F_M.MRAM\[772\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_117_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_1019 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7295__A2 _3606_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7246_ _3294_ _3464_ _3296_ _3584_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
X_4458_ _1126_ _1130_ _1131_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__6342__I1 _2016_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7177_ mod.Data_Mem.F_M.MRAM\[22\]\[3\] _3544_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4389_ mod.Arithmetic.CN.I_in\[28\] _1062_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_98_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6128_ _2695_ _2704_ _2744_ _0064_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_100_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3105 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3116 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6059_ mod.Data_Mem.F_M.MRAM\[14\]\[7\] mod.Data_Mem.F_M.MRAM\[15\]\[7\] _2295_ _2677_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_3127 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_1090 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3138 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2404 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3149 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2415 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2426 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2437 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_148_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2448 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2459 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1714 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_971 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1725 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6558__A1 _2353_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_1017 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6558__B2 _2642_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1736 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1747 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1769 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3947__I _0624_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_154_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_1200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5533__A2 _1729_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_107_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5297__A1 mod.Data_Mem.F_M.MRAM\[783\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7890__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6993__I _3434_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xtiny_user_project_20 io_oeb[9] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_77_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtiny_user_project_31 io_oeb[20] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_77_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtiny_user_project_42 io_oeb[31] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_53 io_out[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_64 io_out[15] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XANTENNA__5049__A1 _1715_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_607 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xtiny_user_project_75 io_out[34] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XANTENNA__6246__B1 _1664_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xtiny_user_project_86 la_data_out[7] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_92_713 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtiny_user_project_97 la_data_out[18] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XANTENNA__8246__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6341__S0 _2448_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5402__I _2062_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4018__I mod.Arithmetic.CN.I_in\[22\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6549__A1 _1966_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2960 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_72_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2971 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_17_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2982 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2993 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_643 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8396__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5072__I1 mod.Data_Mem.F_M.MRAM\[2\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7349__I0 _3620_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_890 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5430_ _2084_ _2085_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5524__A2 _2087_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5361_ mod.Data_Mem.F_M.MRAM\[15\]\[7\] _1886_ _2023_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_58_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__7064__I mod.Data_Mem.F_M.MRAM\[20\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4312_ _0984_ _0985_ _0986_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_7100_ mod.Data_Mem.F_M.MRAM\[23\]\[5\] _3497_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_8080_ _0280_ net1 mod.Data_Mem.F_M.MRAM\[23\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_82_1208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5292_ _1875_ mod.Data_Mem.F_M.MRAM\[768\]\[5\] _1956_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_113_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_7031_ _3459_ _0253_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_102_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4243_ _0842_ _0917_ _0918_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_68_710 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5383__S1 _1590_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4174_ _0825_ _0836_ _0849_ _0850_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_56_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6408__I _2385_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5835__I0 mod.Data_Mem.F_M.MRAM\[14\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_746 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7933_ _0159_ net1 mod.Data_Mem.F_M.MRAM\[8\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_64_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5460__A1 _2069_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7864_ _0090_ net1 mod.Data_Mem.F_M.MRAM\[11\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_23_312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_169_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6815_ _3326_ _0170_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_51_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7795_ _3806_ mod.Data_Mem.F_M.MRAM\[798\]\[5\] _3894_ _3896_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__4015__A2 _0691_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_1001 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6746_ _3249_ mod.Data_Mem.F_M.MRAM\[0\]\[4\] _3279_ _3280_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_3958_ _0634_ _0635_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_104_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_91_1083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6677_ mod.Data_Mem.F_M.dest\[1\] mod.Data_Mem.F_M.dest\[0\] _3231_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_52_1078 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6012__I0 mod.Data_Mem.F_M.MRAM\[16\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_164_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_8416_ _0512_ net1 mod.Data_Mem.F_M.MRAM\[790\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__5515__A2 _2154_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5628_ _2089_ _2099_ _2257_ _2260_ _2261_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_136_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8119__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_105_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8347_ _0443_ net1 mod.Data_Mem.F_M.MRAM\[780\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5559_ _2196_ _2197_ _2198_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_117_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_160_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8278_ _0374_ net1 mod.Data_Mem.F_M.MRAM\[770\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_132_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7229_ _3523_ mod.Data_Mem.F_M.MRAM\[30\]\[0\] _3574_ _3575_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__8269__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5374__S1 _1642_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_58_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_1185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_927 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_150_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_584 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2201 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2212 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2223 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2234 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_162_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_2245 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1500 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2256 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1511 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2267 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1522 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2278 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_40 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_54_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1533 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_51 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_54_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1544 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2289 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_62 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1555 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_14_356 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1566 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5203__A1 _1631_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_148_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_84 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_42_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1577 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_95 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1588 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_35_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_167_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_759 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_584 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5506__A2 mod.Data_Mem.F_M.MRAM\[799\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_155_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_1052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4190__A1 _0863_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_1085 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_604 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_150_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_37_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_116_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7612__I _3797_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5333__S _1892_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_49_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_65_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5132__I _1669_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4245__A2 _0914_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6490__I0 mod.Data_Mem.F_M.MRAM\[12\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4971__I _1600_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4930_ _1598_ _1599_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_45_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5993__A2 mod.Data_Mem.F_M.MRAM\[789\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_166_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_2790 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_127_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4861_ _1529_ _1530_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6600_ _3190_ _0091_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_61_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7580_ _3311_ _3778_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4792_ _0696_ _1460_ _1461_ _1462_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_159_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_20_348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6898__I mod.Data_Mem.F_M.dest\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6531_ _3106_ mod.Data_Mem.F_M.MRAM\[13\]\[6\] _2394_ _3133_ _3134_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_146_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6462_ _3067_ _3068_ _3069_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_118_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8201_ _0086_ net2 net1 mod.I_addr\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_5413_ _2071_ _2072_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6393_ _2866_ _3002_ _0071_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_133_217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5899__I3 mod.Data_Mem.F_M.MRAM\[21\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5344_ _1872_ _2006_ _1884_ _2007_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__8411__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8132_ mod.Data_Mem.F_M.out_data\[42\] net2 net1 mod.Arithmetic.CN.I_in\[42\] vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_142_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_1196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8063_ _0272_ net1 mod.Data_Mem.F_M.MRAM\[21\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5275_ _1931_ _1936_ _1938_ _1563_ _1939_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_99_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_141_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7014_ _3447_ _3448_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_4226_ _0890_ _0900_ _0901_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_102_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4484__A2 _1141_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8561__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4157_ _0655_ mod.Arithmetic.CN.I_in\[40\] mod.Arithmetic.CN.I_in\[41\] _0833_ vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_56_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4088_ _0748_ _0763_ _0764_ _0661_ _0765_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_83_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5433__A1 _2085_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7916_ _0142_ net1 mod.Data_Mem.F_M.MRAM\[10\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_37_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_145_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7847_ mod.Data_Mem.F_M.MRAM\[9\]\[2\] _3926_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_54_1107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_462 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7778_ _3782_ mod.Data_Mem.F_M.MRAM\[797\]\[6\] _3883_ _3886_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_149_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6729_ mod.Data_Mem.F_M.MRAM\[10\]\[7\] _3268_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_20_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_165_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_137_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5217__I _1530_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8091__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4172__A1 _0662_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_965 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3960__I _0636_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5153__S _1816_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5347__S1 _2009_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5672__A1 _2301_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_47_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6492__B _2103_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_1078 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2020 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2031 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_610 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2042 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2053 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2064 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1330 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3986__A1 _0640_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2075 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1341 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2086 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1352 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2097 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_985 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1363 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1374 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1385 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1396 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8434__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8584__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_96_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5060_ _1631_ _1671_ _1727_ _1728_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_42_1000 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_819 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4011_ _0687_ mod.Arithmetic.I_out\[74\] _0684_ mod.Arithmetic.I_out\[73\] _0688_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_2
XANTENNA__5663__A1 _2135_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_713 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_532 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5962_ _2264_ mod.Data_Mem.F_M.MRAM\[20\]\[5\] _2582_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_92_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4769__A3 mod.Arithmetic.CN.I_in\[61\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7701_ _3844_ _0538_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4913_ mod.Data_Mem.F_M.MRAM\[771\]\[0\] mod.Data_Mem.F_M.MRAM\[770\]\[0\] _1581_
+ _1582_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_5893_ _2275_ mod.Data_Mem.F_M.MRAM\[773\]\[3\] _2515_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_7632_ mod.Data_Mem.F_M.MRAM\[788\]\[0\] _3810_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_21_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5718__A2 mod.Data_Mem.F_M.MRAM\[29\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4844_ _1512_ _1513_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_14_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_7563_ _3754_ mod.Data_Mem.F_M.MRAM\[784\]\[5\] _3760_ _3768_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4775_ _1300_ _1321_ _1445_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_147_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6514_ _2475_ _1971_ _2406_ _3117_ _3118_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_7494_ _3724_ _0451_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_119_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_49_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6445_ _3041_ _3052_ _3053_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__7191__I1 mod.Data_Mem.F_M.MRAM\[29\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6376_ _2891_ _2042_ _2986_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_88_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8115_ mod.Data_Mem.F_M.out_data\[25\] net2 net1 mod.Arithmetic.CN.I_in\[25\] vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_5327_ mod.Data_Mem.F_M.MRAM\[3\]\[6\] mod.Data_Mem.F_M.MRAM\[2\]\[6\] _1877_ _1990_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_88_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_646 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7951__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8046_ _0255_ net1 mod.Data_Mem.F_M.MRAM\[18\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_76_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5258_ _1704_ _1922_ _1923_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_102_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5654__A1 _2068_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_1144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4209_ mod.Arithmetic.CN.I_in\[8\] _0707_ _0814_ _0883_ _0884_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
X_5189_ mod.Data_Mem.F_M.MRAM\[768\]\[3\] _1855_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_112_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_830 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_746 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_1188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8307__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5257__I1 mod.Data_Mem.F_M.MRAM\[784\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_429 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5500__I _2059_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5957__A2 _2555_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_1062 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__8457__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5709__A2 mod.Data_Mem.F_M.MRAM\[28\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_169_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_106_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4768__I0 mod.Arithmetic.ACTI.x\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6221__I3 mod.Data_Mem.F_M.MRAM\[4\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3955__I _0613_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6382__A2 _2990_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4393__A1 _0642_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4145__A1 _0621_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_1191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5893__A1 _2275_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_152_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_105_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_78_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_819 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5645__A1 _2270_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6506__I _2107_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5948__A2 mod.Data_Mem.F_M.MRAM\[3\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5410__I _1595_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4026__I _0702_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1160 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1171 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_63_81 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_1195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1182 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6748__I1 mod.Data_Mem.F_M.MRAM\[0\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1193 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_169_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7570__A1 _3705_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6373__A2 _2041_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4560_ _1226_ _1231_ _1232_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_156_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4491_ _1075_ _1076_ _1163_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__6125__A2 _1497_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4136__A1 _0639_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7974__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6230_ _2831_ _2834_ _2835_ _2093_ _2843_ _2844_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_98_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_1111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6161_ _2681_ _2772_ _2776_ _2777_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_83_1144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_911 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_83_1155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_933 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5112_ _1579_ _1779_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6092_ _1764_ _1613_ _2709_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_83_1199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_465 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_966 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5636__A1 _2266_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4439__A2 mod.Arithmetic.CN.I_in\[57\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_977 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6684__I0 _3228_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_988 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5043_ _1707_ mod.Data_Mem.F_M.MRAM\[771\]\[1\] _1710_ _1711_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_80_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6994_ _3386_ mod.Data_Mem.F_M.MRAM\[17\]\[0\] _3435_ _3436_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_80_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6987__I1 mod.Data_Mem.F_M.MRAM\[16\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6061__A1 _2410_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5945_ _1533_ _2137_ _2557_ _2564_ _2565_ _2566_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_90_1104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5876_ _2496_ _2497_ _2378_ _2498_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_21_432 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7615_ _3747_ mod.Data_Mem.F_M.MRAM\[787\]\[1\] _3798_ _3800_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4827_ _1494_ _1495_ _1496_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_8595_ _0611_ net1 mod.Instr_Mem.instruction\[30\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__7247__I _3584_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4375__A1 _0968_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5195__C _1490_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7546_ _3731_ mod.Data_Mem.F_M.MRAM\[783\]\[7\] _3752_ _3757_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4758_ _1421_ _1427_ _1428_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_119_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_146_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7477_ _3714_ _0444_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4689_ _1225_ _1354_ _0997_ _1360_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__4127__A1 _0633_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_1066 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6428_ _1933_ mod.Data_Mem.F_M.MRAM\[769\]\[1\] _3036_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_162_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_88_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6359_ mod.Data_Mem.F_M.MRAM\[781\]\[6\] _2751_ _2902_ mod.Data_Mem.F_M.MRAM\[780\]\[6\]
+ _2969_ _2970_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_68_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_89_977 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_765 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5627__A1 _2258_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5478__I1 mod.Data_Mem.F_M.MRAM\[799\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8029_ _0238_ net1 mod.Data_Mem.F_M.MRAM\[16\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_29_532 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_75_148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6052__A1 _2539_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_568 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4063__B1 _0703_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_210 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_13_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_24_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_254 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_287 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_8_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_33_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7997__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_166_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_149_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_138_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_165_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_158_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5866__A1 _2447_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4669__A2 _1339_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5618__A1 mod.Data_Mem.F_M.MRAM\[29\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5618__B2 mod.Data_Mem.F_M.MRAM\[28\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_584 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5341__S _1906_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6830__A3 _3335_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_682 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6043__A1 _2434_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3991_ _0660_ _0667_ _0668_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_5730_ _2354_ _2355_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_31_752 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5661_ _2287_ _2289_ _2291_ _2292_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_88_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7400_ _3673_ _0408_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__8002__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4612_ _1165_ _1187_ _1283_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_8380_ _0476_ net1 mod.Data_Mem.F_M.MRAM\[784\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5592_ _1811_ _2229_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_157_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7331_ _3603_ mod.Data_Mem.F_M.MRAM\[771\]\[0\] _3636_ _3637_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4543_ mod.Arithmetic.CN.I_in\[35\] _1091_ _1215_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_11_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_85_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7262_ _3593_ _0350_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4474_ _1035_ _1036_ _1145_ _1147_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_144_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__8152__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5857__A1 _2383_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6213_ _2824_ _2825_ _2826_ _2827_ _2686_ _2828_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
X_7193_ _3549_ _3553_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_48_1083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_540 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6144_ _2360_ mod.Data_Mem.F_M.MRAM\[6\]\[1\] mod.Data_Mem.F_M.MRAM\[7\]\[1\] _2188_
+ _2760_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_730 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_903 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_752 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5609__A1 _1953_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_785 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6075_ _2691_ _2692_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_796 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5026_ _1691_ mod.Data_Mem.F_M.MRAM\[791\]\[1\] _1693_ _1694_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_2608 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_66_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_513 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2619 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_546 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6034__A1 _2549_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1907 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1918 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_568 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1929 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6977_ _3425_ _0233_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_80_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7782__A1 _3294_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_1010 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5928_ _2144_ _2549_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_55_1032 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_730 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_1122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_142_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6337__A2 _2003_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_1087 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5859_ _2435_ _2477_ _2478_ _2439_ _2481_ _2482_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_148_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_8578_ _0594_ net1 mod.Instr_Mem.instruction\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_21_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7529_ _3746_ _0464_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_5_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_147_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7137__I1 mod.Data_Mem.F_M.MRAM\[19\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_163_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5848__A1 _2428_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_730 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_752 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4520__A1 mod.Arithmetic.CN.I_in\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtiny_user_project_104 la_data_out[25] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_0_177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_103_584 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xtiny_user_project_115 la_data_out[36] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_62_1069 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5161__S _1685_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xtiny_user_project_126 la_data_out[47] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_137 la_data_out[58] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_148 wbs_dat_o[1] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_76_468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtiny_user_project_159 wbs_dat_o[12] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_91_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5895__I _2116_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_836 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8025__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_160_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_9_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_157_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_1198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5000__A2 _1667_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8175__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7128__I1 mod.Data_Mem.F_M.MRAM\[19\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_158_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_126_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6500__A2 mod.Data_Mem.F_M.MRAM\[768\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7551__S _3760_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_1059 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4190_ _0863_ _0864_ _0865_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_79_251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_1125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7300__I1 mod.Data_Mem.F_M.MRAM\[768\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6264__A1 _2876_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_800 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_48_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4814__A2 _1483_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6900_ _3373_ _3374_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_78_1010 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7880_ _0106_ net1 mod.Data_Mem.F_M.MRAM\[26\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_63_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6016__A1 _1685_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6831_ _3336_ _3337_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_63_674 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6567__A2 _3158_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4923__B _1558_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6762_ mod.Data_Mem.F_M.MRAM\[8\]\[4\] _3288_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_3974_ _0650_ _0651_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_52_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_8501_ _0005_ net1 mod.Data_Mem.F_M.out_data\[77\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5713_ _2339_ mod.Data_Mem.F_M.MRAM\[796\]\[6\] _2311_ _2340_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__8518__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6693_ _3244_ _0130_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6319__A2 _1937_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5790__A3 _2374_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8432_ _0528_ net1 mod.Data_Mem.F_M.MRAM\[792\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__5378__I0 mod.Data_Mem.F_M.MRAM\[769\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5644_ _2275_ mod.Data_Mem.F_M.MRAM\[796\]\[1\] _2268_ _2276_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_15_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_163_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_8363_ _0459_ net1 mod.Data_Mem.F_M.MRAM\[782\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_129_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5575_ mod.Data_Mem.F_M.MRAM\[29\]\[3\] _2213_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_102_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_1161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7314_ _3610_ _3626_ _3627_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__7819__A2 mod.I_addr\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4526_ _1103_ _1198_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_117_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8294_ _0390_ net1 mod.Data_Mem.F_M.MRAM\[772\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_132_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_145_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_7245_ _3583_ _0343_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_85_1058 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4457_ _1127_ _1129_ _1130_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_104_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4502__A1 _0613_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7176_ _3543_ _0314_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_58_402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4388_ _0632_ _1061_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_86_711 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6127_ _1726_ _2727_ _2735_ _2742_ _2743_ _2744_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XTAP_571 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3106 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_46_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6058_ _2062_ mod.Data_Mem.F_M.MRAM\[5\]\[7\] _2675_ _2572_ _2676_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_86_788 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3117 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_61_1080 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3128 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3139 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_682 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2405 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5009_ _1676_ _1677_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__8048__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2416 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2427 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2438 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2449 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1704 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1715 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_983 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_1007 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_1127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1726 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6558__A2 _2347_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1737 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_121_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_1149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1748 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4569__A1 _0614_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_858 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1759 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5766__B1 _2390_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8198__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7507__A1 _3634_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_891 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_155_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3963__I _0613_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_1212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_151_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5297__A2 _1599_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_819 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_110_307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6495__B _3099_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtiny_user_project_21 io_oeb[10] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_32 io_oeb[21] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_1_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xtiny_user_project_43 io_oeb[32] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_54 io_out[5] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_65 io_out[24] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_77_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtiny_user_project_76 io_out[35] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_77_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xtiny_user_project_87 la_data_out[8] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_98 la_data_out[19] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_18_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6341__S1 _1932_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7046__I0 _3452_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_972 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_1216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2950 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2961 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8227__RN net2 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2972 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2983 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2994 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7349__I1 mod.Data_Mem.F_M.MRAM\[771\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7546__S _3752_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4034__I mod.Arithmetic.I_out\[73\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_145_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_126_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5360_ _2022_ _0006_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_114_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_126_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4311_ _0897_ _0833_ _0896_ mod.Arithmetic.CN.I_in\[41\] _0985_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_141_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5291_ mod.Data_Mem.F_M.MRAM\[769\]\[5\] _1955_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__6485__A1 _2072_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7030_ _3416_ mod.Data_Mem.F_M.MRAM\[18\]\[5\] _3457_ _3459_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4242_ _0615_ mod.Arithmetic.ACTI.x\[2\] _0917_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_45_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_1053 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4173_ _0837_ _0839_ _0848_ _0849_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XANTENNA__7080__I mod.Data_Mem.F_M.MRAM\[21\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6237__A1 _1931_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7285__I0 _3603_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5835__I1 mod.Data_Mem.F_M.MRAM\[15\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_82_213 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7932_ _0158_ net1 mod.Data_Mem.F_M.MRAM\[8\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_83_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7863_ _0089_ net1 mod.Data_Mem.F_M.MRAM\[11\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_82_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8340__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_611 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6814_ mod.Data_Mem.F_M.MRAM\[789\]\[2\] _3326_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_51_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7794_ _3895_ _0580_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__7908__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_168_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6745_ _3273_ _3279_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_11_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_1051 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_1013 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3957_ _0633_ _0634_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_91_1062 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8490__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6676_ _3229_ _3230_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_52_1068 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6012__I1 mod.Data_Mem.F_M.MRAM\[17\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8498__D _0002_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8415_ _0511_ net1 mod.Data_Mem.F_M.MRAM\[788\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5627_ _2258_ mod.Data_Mem.F_M.MRAM\[796\]\[0\] _2259_ _2260_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_136_237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_118_974 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4723__A1 _1031_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8346_ _0442_ net1 mod.Data_Mem.F_M.MRAM\[780\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5558_ _2189_ mod.Data_Mem.F_M.MRAM\[799\]\[2\] mod.Data_Mem.F_M.MRAM\[798\]\[2\]
+ _1915_ _2197_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_133_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_933 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4509_ _1177_ _1179_ _1175_ _1181_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_8277_ _0373_ net1 mod.Data_Mem.F_M.MRAM\[770\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__7191__S _3550_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5489_ _2059_ _2134_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_132_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6476__A1 _2184_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_988 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7228_ _3573_ _3574_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_59_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_1153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7159_ _3248_ _3533_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_58_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_47_906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6228__A1 mod.Data_Mem.F_M.MRAM\[13\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_390 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_59_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_1197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_46_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2202 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5987__B1 _2606_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2213 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2224 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7028__I0 _3456_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2235 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2246 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1501 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1512 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2257 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3958__I _0634_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_30 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_70_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2268 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1523 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_931 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2279 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_41 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_15_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1534 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_155_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_52 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1545 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_63 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1556 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1036 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_74 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1567 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_85 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1578 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1058 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_96 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_70_997 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1589 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6270__S _1742_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5394__B _2055_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6164__B1 _1703_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7165__I _3255_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_157_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_109_974 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_109_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_108_473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_68_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8213__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6467__A1 _2171_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_817 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_155_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_124_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_81_1220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5413__I _2071_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6219__A1 _2567_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8363__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_972 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6490__I1 mod.Data_Mem.F_M.MRAM\[14\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_983 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_1002 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_1182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2780 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_430 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4860_ _1501_ _1528_ _1529_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_2791 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4791_ mod.Arithmetic.CN.I_in\[23\] mod.Arithmetic.CN.I_in\[31\] _1461_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_20_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6530_ _2424_ mod.Data_Mem.F_M.MRAM\[12\]\[6\] _3133_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_119_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_6461_ mod.Data_Mem.F_M.MRAM\[12\]\[2\] _1886_ _2536_ _2486_ _3068_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_8200_ _0085_ net2 net1 mod.I_addr\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_51_1090 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4705__A1 _0632_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5412_ _2070_ _2071_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6392_ _2868_ _2993_ _3001_ _3002_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_115_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8131_ mod.Data_Mem.F_M.out_data\[41\] net2 net1 mod.Arithmetic.CN.I_in\[41\] vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_5343_ _2002_ _2003_ _2004_ _2005_ _1910_ _1590_ _2006_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_115_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_47_1126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_114_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6458__A1 _2063_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8062_ _0271_ net1 mod.Data_Mem.F_M.MRAM\[20\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_82_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5274_ _1645_ _1937_ _1938_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_102_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7013_ _3433_ _3446_ _3421_ _3447_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_4225_ _0895_ _0899_ _0900_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__5130__A1 mod.Data_Mem.F_M.MRAM\[799\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4156_ _0657_ _0831_ _0832_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_95_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_96_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4087_ _0706_ _0751_ _0745_ _0764_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XANTENNA__5433__A2 _2087_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7915_ _0141_ net1 mod.Data_Mem.F_M.MRAM\[10\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_36_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__4383__B _0809_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_1124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_169_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7846_ _3925_ _0601_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_19_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_1157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_975 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7880__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7777_ _3885_ _0573_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4989_ _1655_ _1656_ _1657_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_51_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6728_ _3267_ _0142_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_109_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6659_ mod.Data_Mem.F_M.MRAM\[27\]\[1\] _3220_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__8236__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_152_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8329_ _0425_ net1 mod.Data_Mem.F_M.MRAM\[777\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_79_806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7497__I0 _3725_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6449__A1 _3017_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__8386__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5121__A1 _1715_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5233__I _1799_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_1062 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_574 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_46_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2010 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_62_717 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_74_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2021 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2032 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2043 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5975__A3 _2594_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2054 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1320 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2065 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1331 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3986__A2 mod.Arithmetic.CN.I_in\[64\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2076 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1342 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_1208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2087 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1353 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2098 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1364 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1375 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5188__A1 _1745_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_159_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1397 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_161_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_156_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6137__B1 mod.Data_Mem.F_M.MRAM\[15\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5408__I _2068_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_155_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4163__A2 _0838_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5143__I _1543_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_1050 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4010_ _0682_ _0687_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XANTENNA__5663__A2 mod.Data_Mem.F_M.MRAM\[29\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_503 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_18_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5961_ _2475_ mod.Data_Mem.F_M.MRAM\[21\]\[5\] _2581_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_80_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8109__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4769__A4 _1366_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7700_ mod.Data_Mem.F_M.MRAM\[793\]\[2\] _3844_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_80_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4912_ _1580_ _1581_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__6903__S _3376_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_430 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5892_ _2511_ _1851_ _2513_ _2514_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_7631_ _2049_ _3804_ _3809_ _0503_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_61_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4843_ _1502_ _1512_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_33_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8259__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7562_ _3767_ _0476_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4774_ _1435_ _1438_ _1443_ _1444_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
X_6513_ _2528_ mod.Data_Mem.F_M.MRAM\[0\]\[5\] _3117_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_146_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_20_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_119_546 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7493_ _3711_ mod.Data_Mem.F_M.MRAM\[781\]\[3\] _3720_ _3724_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_88_1204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_1106 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4222__I mod.Arithmetic.CN.I_in\[42\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6444_ _3045_ _3048_ _3051_ _2831_ _2073_ _3052_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_134_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_538 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5351__A1 _1903_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4154__A2 _0829_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6375_ _2779_ _2983_ _2984_ _2985_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_161_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7533__I _3305_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8114_ mod.Data_Mem.F_M.out_data\[24\] net2 net1 mod.Arithmetic.CN.I_in\[24\] vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_5326_ mod.Data_Mem.F_M.MRAM\[1\]\[6\] mod.Data_Mem.F_M.MRAM\[0\]\[6\] _1609_ _1989_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_103_914 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_103_936 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6149__I _2706_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8045_ _0254_ net1 mod.Data_Mem.F_M.MRAM\[18\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_130_755 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5257_ mod.Data_Mem.F_M.MRAM\[785\]\[4\] mod.Data_Mem.F_M.MRAM\[784\]\[4\] _1580_
+ _1922_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_87_146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5654__A2 _2285_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4208_ mod.Arithmetic.CN.I_in\[8\] _0814_ _0882_ _0883_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_75_319 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_894 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5188_ _1745_ _1853_ _1854_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_60_1156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4139_ _0631_ _0814_ _0815_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_44_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4209__A3 _0814_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_503 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_897 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_249 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7829_ _3174_ _3909_ _3908_ _3915_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_169_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_1017 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_138_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_31 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_165_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_137_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_153_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4145__A2 _0656_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6390__I0 _2252_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5164__S _1829_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_603 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5893__A2 mod.Data_Mem.F_M.MRAM\[773\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_156_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_3_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5645__A2 _2122_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_94_639 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_35_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_897 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_867 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_878 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8401__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_1163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1161 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1172 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4751__B _1340_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5339__S _1814_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1183 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1194 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4908__A1 _1563_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7570__A2 _3335_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_128_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5138__I _1799_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8551__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4490_ _1160_ _1082_ _1161_ _1162_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_6_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6381__I0 _2051_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7353__I mod.Data_Mem.F_M.MRAM\[772\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6160_ _1661_ _2773_ _2774_ _2775_ _2776_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_135_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_901 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_124_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_923 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_69_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5111_ _1690_ _1778_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_83_1167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_755 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_945 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6091_ _2707_ _2708_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_978 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4439__A3 _0922_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5042_ _1708_ _1709_ _1710_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_38_500 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_820 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6993_ _3434_ _3435_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_19_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__8081__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5944_ _2065_ _2565_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_34_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_168_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5875_ mod.Data_Mem.F_M.MRAM\[786\]\[3\] mod.Data_Mem.F_M.MRAM\[787\]\[3\] _1932_
+ _2497_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_7614_ _3799_ _0496_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4826_ mod.Data_Mem.F_M.src\[4\] _1495_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_8594_ _0610_ net1 mod.Instr_Mem.instruction\[24\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_7545_ _3756_ _0470_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4375__A2 _0965_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_147_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_21_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4757_ _1422_ _1426_ _1427_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_119_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7476_ _3615_ mod.Data_Mem.F_M.MRAM\[780\]\[4\] _3713_ _3714_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4688_ _1353_ _1357_ _1358_ _1359_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__4127__A2 mod.Arithmetic.CN.I_in\[17\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6427_ _2728_ mod.Data_Mem.F_M.MRAM\[781\]\[1\] _2381_ _3034_ _3035_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_135_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_1029 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6358_ _2752_ _2968_ _2969_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_88_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5309_ _1769_ _1971_ _1972_ _1973_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_130_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6289_ _1543_ _2902_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_8028_ _0237_ net1 mod.Data_Mem.F_M.MRAM\[16\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_75_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_76_639 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__8424__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_72_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6052__A2 _2663_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_1049 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4063__B2 mod.Arithmetic.CN.I_in\[22\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_31_219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_233 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__8574__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3966__I _0642_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_255 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_8519__183 net183 vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_24_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_277 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_129_107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5938__I0 mod.Data_Mem.F_M.MRAM\[16\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_288 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_126_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_165_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_79_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6115__I0 mod.Data_Mem.F_M.MRAM\[7\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5618__A2 _2086_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_871 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_893 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_58_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_75_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5421__I _2078_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7615__I0 _3747_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_1214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_171 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_165_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6043__A2 _2660_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_165_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3990_ _0662_ _0666_ _0667_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_50_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5660_ _2290_ _2125_ _2291_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__7941__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4611_ _1197_ _1280_ _1281_ _1282_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__5554__A1 _2184_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_30_285 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5591_ _1606_ _2228_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_7330_ _3635_ _3636_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_8_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_102_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4542_ _0636_ mod.Arithmetic.CN.I_in\[36\] _0892_ _0980_ _1214_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
X_7261_ mod.Data_Mem.F_M.MRAM\[31\]\[6\] _3319_ _3590_ _3593_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_116_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4473_ _1035_ _1036_ _1145_ _1146_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or3_1
X_6212_ _1734_ _1789_ _2775_ _2827_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__5857__A2 mod.Data_Mem.F_M.MRAM\[773\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7192_ _3552_ _0321_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_98_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6143_ _2691_ _2759_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_48_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8447__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_753 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5609__A2 mod.Data_Mem.F_M.MRAM\[31\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_714 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6074_ _2685_ _2691_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_797 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_1213 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5025_ _1692_ mod.Data_Mem.F_M.MRAM\[790\]\[1\] _1693_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_100_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4293__A1 _0878_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2609 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_66_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1908 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1919 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6976_ _3393_ mod.Data_Mem.F_M.MRAM\[16\]\[1\] _3423_ _3425_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__5093__I0 _1755_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_675 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_1180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5927_ _2396_ _2548_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_94_1082 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5858_ _2440_ _2479_ _2480_ _2481_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_4809_ _1372_ _1380_ _1478_ _1479_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__7194__S _3553_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8577_ _0593_ net1 mod.Instr_Mem.instruction\[26\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5789_ _2413_ _2414_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_108_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7528_ _3718_ mod.Data_Mem.F_M.MRAM\[783\]\[0\] _3745_ _3746_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_107_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7459_ mod.Data_Mem.F_M.MRAM\[778\]\[6\] _3703_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_107_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_162_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_107_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_1184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_103_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtiny_user_project_105 la_data_out[26] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_116 la_data_out[37] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_76_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtiny_user_project_127 la_data_out[48] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_138 la_data_out[59] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_64_609 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xtiny_user_project_149 wbs_dat_o[2] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_91_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_642 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7964__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7168__I _3258_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_1133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6072__I _2681_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_1155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_40_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_94 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_154_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_5_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_153_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_81 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_872 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_140_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_132_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_95_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_1159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_745 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_393 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6264__A2 _1878_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5311__I1 _1970_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_82_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_1033 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6016__A2 mod.Data_Mem.F_M.MRAM\[19\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4990__I _1646_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6830_ _3332_ _3298_ _3335_ _3336_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_36_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_23_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_984 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_1200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6761_ _3287_ _0155_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_62_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5775__A1 _2313_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_859 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3973_ _0645_ _0650_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_5712_ _2025_ _2339_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_50_358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8500_ _0004_ net1 mod.Data_Mem.F_M.out_data\[76\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6692_ _3243_ mod.Data_Mem.F_M.MRAM\[28\]\[2\] _3237_ _3244_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_8431_ _0527_ net1 mod.Data_Mem.F_M.MRAM\[791\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5643_ _1586_ _2275_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__5378__I1 mod.Data_Mem.F_M.MRAM\[768\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8362_ _0458_ net1 mod.Data_Mem.F_M.MRAM\[782\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_157_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5574_ _1601_ _2212_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_102_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7313_ _3625_ _3626_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4525_ _1159_ _1162_ _1196_ _1197_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
X_8293_ _0389_ net1 mod.Data_Mem.F_M.MRAM\[772\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_89_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_102_1086 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_1037 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7244_ _3539_ mod.Data_Mem.F_M.MRAM\[30\]\[7\] _3579_ _3583_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_116_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4456_ _1008_ _1128_ _1129_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_137_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_131_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7175_ mod.Data_Mem.F_M.MRAM\[22\]\[2\] _3543_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_59_904 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4387_ _0956_ _1059_ _1060_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6126_ _2366_ _2195_ _2743_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XTAP_561 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_572 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6057_ _2288_ mod.Data_Mem.F_M.MRAM\[4\]\[7\] _2675_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XTAP_3107 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4266__A1 _0768_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5061__I _1728_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3118 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3129 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7987__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5008_ _1593_ _1676_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_96_1111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2406 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2417 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2428 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7189__S _3550_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2439 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_148_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1705 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1716 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1727 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1749 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5766__A1 _2388_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4569__A2 mod.Arithmetic.CN.I_in\[69\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6959_ _3413_ _0227_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_53_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5766__B2 _2290_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7995__RN net2 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8516__186 net186 vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_139_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_136_942 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_163_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_100_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_107_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_135_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8172__RN net2 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_151_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xtiny_user_project_11 io_oeb[0] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_104_872 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6495__C _2108_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xtiny_user_project_22 io_oeb[11] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XANTENNA__5129__S0 _1527_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_680 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xtiny_user_project_33 io_oeb[22] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_49_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtiny_user_project_44 io_oeb[33] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_103_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xtiny_user_project_55 io_out[6] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_103_393 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtiny_user_project_66 io_out[25] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XANTENNA__6246__A2 _2221_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xtiny_user_project_77 io_out[36] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_64_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xtiny_user_project_88 la_data_out[9] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XANTENNA__4257__A1 _0824_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xtiny_user_project_99 la_data_out[20] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_58_981 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_322 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7046__I1 mod.Data_Mem.F_M.MRAM\[1\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2940 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_17_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2951 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2962 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2973 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_32_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2984 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8142__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2995 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7986__RN net2 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_678 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_41_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8292__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6182__A1 _2073_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_161_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6309__I0 _1978_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5146__I _1811_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4310_ _0983_ _0984_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_5290_ _1953_ _1954_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_99_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4241_ _0915_ mod.Arithmetic.ACTI.x\[1\] _0663_ _0916_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__6485__A2 _2509_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8163__RN net2 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_68_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4172_ _0662_ _0841_ _0847_ _0848_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_67_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7285__I1 mod.Data_Mem.F_M.MRAM\[768\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6237__A2 _1848_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_575 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_981 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7931_ _0157_ net1 mod.Data_Mem.F_M.MRAM\[8\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__5996__A1 _2313_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4799__A2 _1176_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7862_ _0088_ net1 mod.Data_Mem.F_M.MRAM\[11\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_35_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_461 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6813_ _3325_ _0169_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5748__A1 _1542_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6796__I0 mod.Data_Mem.F_M.MRAM\[799\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7793_ _3312_ mod.Data_Mem.F_M.MRAM\[798\]\[4\] _3894_ _3895_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_50_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_1161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6744_ _3278_ _0147_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_3956_ _0632_ _0633_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4420__A1 _0828_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_1025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6675_ mod.Data_Mem.F_M.dest\[4\] mod.Data_Mem.F_M.dest\[2\] _3229_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__5257__S _1580_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8414_ _0510_ net1 mod.Data_Mem.F_M.MRAM\[788\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5626_ _2216_ _2259_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_8345_ _0441_ net1 mod.Data_Mem.F_M.MRAM\[780\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5557_ _1644_ _2196_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_117_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5056__I mod.Data_Mem.F_M.src\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_151_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_145_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_132_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4508_ _1175_ _1177_ _1179_ _1180_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or3_1
X_8276_ _0372_ net1 mod.Data_Mem.F_M.MRAM\[770\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_117_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5488_ _2114_ _2128_ _2131_ _2133_ _0035_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_133_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4895__I _1525_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6476__A2 _3079_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7227_ _3230_ _3464_ _3389_ _3573_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__8154__RN net2 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4439_ _0650_ mod.Arithmetic.CN.I_in\[57\] _0922_ _1019_ _1112_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XANTENNA__7271__I mod.Data_Mem.F_M.MRAM\[5\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8015__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_1132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_150_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_7158_ _3532_ _0307_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_101_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_1165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_380 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6109_ _2692_ _2721_ _2725_ _2726_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__6228__A2 _1729_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_391 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_7089_ _3491_ _0279_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4239__A1 _0615_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_46_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_726 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5987__A1 _2406_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8165__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_759 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2203 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5987__B2 _2403_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2214 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7028__I1 mod.Data_Mem.F_M.MRAM\[18\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2225 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2236 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2247 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1502 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_148_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2258 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_20 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1513 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2269 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_31 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1524 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_42 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_14_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1535 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_81_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1546 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6787__I0 mod.Data_Mem.F_M.MRAM\[799\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_64 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_75 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1568 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_86 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1579 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_148_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_35_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4411__A1 _0988_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3974__I _0650_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_168_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_1158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6164__A1 _1555_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_575 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6164__B2 _1566_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_942 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_143_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_108_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__6467__A2 mod.Data_Mem.F_M.MRAM\[0\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8145__RN net2 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_104_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_391 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8508__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6219__A2 _2572_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5978__A1 _2385_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_951 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6490__I2 mod.Data_Mem.F_M.MRAM\[13\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_1161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_1194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2770 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2781 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2792 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4045__I mod.Arithmetic.CN.I_in\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_162_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4790_ _1307_ _1314_ _1460_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__4402__A1 _1052_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6260__I _2706_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_158_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6460_ _3021_ _2490_ _3066_ _3031_ _3047_ _3067_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_9_362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6155__A1 _1910_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5411_ _2069_ _2070_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_63_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6391_ _2867_ _3000_ _3001_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__4705__A2 mod.Arithmetic.ACTI.x\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_901 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8038__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_8130_ mod.Data_Mem.F_M.out_data\[40\] net2 net1 mod.Arithmetic.CN.I_in\[40\] vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_5342_ mod.Data_Mem.F_M.MRAM\[775\]\[6\] mod.Data_Mem.F_M.MRAM\[774\]\[6\] _1908_
+ _2005_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_86_1154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8061_ _0270_ net1 mod.Data_Mem.F_M.MRAM\[20\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_47_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__8136__RN net2 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_1018 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6458__A2 _3064_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5273_ mod.Data_Mem.F_M.MRAM\[791\]\[5\] mod.Data_Mem.F_M.MRAM\[790\]\[5\] _1783_
+ _1937_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_99_155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7012_ _3388_ _3446_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_4224_ _0896_ _0897_ _0898_ _0899_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__5130__A2 _1775_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8188__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_29_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4155_ _0655_ mod.Arithmetic.CN.I_in\[41\] _0831_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_96_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_575 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4086_ _0749_ _0762_ _0710_ _0763_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__5969__A1 _2588_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7914_ _0140_ net1 mod.Data_Mem.F_M.MRAM\[10\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__5433__A3 _2076_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_1114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_943 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7845_ mod.Data_Mem.F_M.MRAM\[9\]\[1\] _3925_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_168_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_93_1169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_12_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6371__S _2180_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7776_ _3806_ mod.Data_Mem.F_M.MRAM\[797\]\[5\] _3883_ _3885_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4988_ mod.Data_Mem.F_M.MRAM\[17\]\[1\] mod.Data_Mem.F_M.MRAM\[16\]\[1\] _1519_ _1656_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_6727_ mod.Data_Mem.F_M.MRAM\[10\]\[6\] _3267_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_3939_ _0616_ _0617_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6658_ _3219_ _0120_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__7194__I0 _3529_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_249 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5609_ _1953_ mod.Data_Mem.F_M.MRAM\[31\]\[6\] mod.Data_Mem.F_M.MRAM\[30\]\[6\] _2229_
+ _2244_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XANTENNA__6941__I0 _3253_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6589_ _3184_ _0086_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_8328_ _0424_ net1 mod.Data_Mem.F_M.MRAM\[777\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_11_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_1216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8127__RN net2 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7497__I1 mod.Data_Mem.F_M.MRAM\[781\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8259_ _0355_ net1 mod.Data_Mem.F_M.MRAM\[5\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_105_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5121__A2 _1787_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2000 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6082__B1 _2212_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2011 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2022 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_461 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2033 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4632__A1 mod.Arithmetic.CN.I_in\[37\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2044 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1310 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2055 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1321 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2066 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1332 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2077 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_1343 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2088 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1354 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2099 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1365 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_615 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6385__A1 _1565_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1376 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5188__A2 _1853_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1387 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1398 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_126_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_503 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_1023 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6137__A1 _2009_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6137__B2 _1968_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_116_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_569 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6932__I0 _3395_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4699__A1 _0891_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5896__B1 _2516_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8330__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__8118__RN net2 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5424__I _1701_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_111_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_97_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_1084 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8480__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6299__S1 _2759_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5960_ mod.Data_Mem.F_M.MRAM\[16\]\[5\] mod.Data_Mem.F_M.MRAM\[17\]\[5\] _2283_ _2580_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__4623__A1 mod.Arithmetic.CN.I_in\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4911_ _1579_ _1580_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_5891_ _2512_ mod.Data_Mem.F_M.MRAM\[771\]\[3\] _2513_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_7630_ _3322_ _3798_ _3809_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_4842_ mod.Data_Mem.F_M.MRAM\[21\]\[0\] mod.Data_Mem.F_M.MRAM\[20\]\[0\] _1510_ _1511_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__6376__A1 _2891_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_92_1180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7561_ _3725_ mod.Data_Mem.F_M.MRAM\[784\]\[4\] _3760_ _3767_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4773_ _1440_ _1439_ _1442_ _1443_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_105_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6512_ _2696_ mod.Data_Mem.F_M.MRAM\[12\]\[5\] _2596_ _3116_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_7492_ _3723_ _0450_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_88_1216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_162_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6443_ _3049_ _2285_ _3050_ _2453_ _2460_ _2496_ _3051_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_1
X_6374_ _2891_ _2040_ _2984_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_115_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5351__A2 mod.Data_Mem.F_M.MRAM\[786\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7628__A1 _3319_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5325_ mod.Data_Mem.F_M.MRAM\[7\]\[6\] mod.Data_Mem.F_M.MRAM\[6\]\[6\] _1873_ _1988_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_8113_ mod.Data_Mem.F_M.out_data\[23\] net2 net1 mod.Arithmetic.CN.I_in\[23\] vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XANTENNA__8109__RN net2 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_904 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7750__S _3867_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_797 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8044_ _0253_ net1 mod.Data_Mem.F_M.MRAM\[18\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5256_ _1918_ _1919_ _1920_ _1921_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__6300__A1 _2703_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4207_ _0813_ _0715_ _0882_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5187_ _1845_ mod.Data_Mem.F_M.MRAM\[771\]\[3\] _1852_ _1853_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_56_501 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4138_ _0813_ _0709_ _0814_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_60_1168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4069_ _0706_ _0745_ _0746_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_58_1020 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4090__A2 _0708_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8203__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7828_ _3914_ _0595_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6367__A1 _1834_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_924 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_1220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_145_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_51_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7759_ _3782_ mod.Data_Mem.F_M.MRAM\[796\]\[6\] _3872_ _3875_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_156_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_40_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5509__I _2144_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4393__A3 _1062_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__8353__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6914__I0 _3253_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_152_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4145__A3 _0820_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6390__I1 _2255_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_1171 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_3_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_121_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_105_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_101_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_47_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_504 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6803__I _3318_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1140 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1151 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6358__A1 _2752_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1162 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1184 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1195 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_8_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5581__A2 _2179_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_155_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_878 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6905__I0 _3240_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5869__C2 _2170_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6530__A1 _2424_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6381__I1 _2052_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_83_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_913 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5110_ _1759_ _1774_ _1776_ _1508_ _1777_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_124_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_924 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_935 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6090_ _2706_ _2707_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_946 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_83_1179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_69_158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_607 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7870__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4993__I _1639_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_968 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5041_ mod.Data_Mem.F_M.MRAM\[770\]\[1\] _1709_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__4439__A4 _1019_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6914__S _3381_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_504 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8226__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6992_ _3433_ _3371_ _3421_ _3434_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_1213 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6061__A3 _2676_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5943_ _2558_ _2559_ _2563_ _2564_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_40_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6349__A1 _2869_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5874_ _2495_ _2496_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_33_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_167_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7613_ _3771_ mod.Data_Mem.F_M.MRAM\[787\]\[0\] _3798_ _3799_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__8376__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4825_ mod.Data_Mem.F_M.src\[2\] _1494_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_138_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_8593_ _0609_ net1 mod.Instr_Mem.instruction\[17\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__5021__A1 _1685_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7544_ _3729_ mod.Data_Mem.F_M.MRAM\[783\]\[6\] _3752_ _3756_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4756_ mod.Arithmetic.CN.I_in\[39\] _1425_ _1426_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_107_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7475_ _3706_ _3713_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_4687_ _1353_ _1356_ _1358_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_134_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6426_ _2301_ mod.Data_Mem.F_M.MRAM\[780\]\[1\] _3034_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__6521__A1 _2567_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_161_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_150_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6357_ _2904_ mod.Data_Mem.F_M.MRAM\[783\]\[6\] mod.Data_Mem.F_M.MRAM\[782\]\[6\]
+ _2905_ _2968_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_103_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5308_ _1942_ mod.Data_Mem.F_M.MRAM\[0\]\[5\] _1972_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_62_1208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_130_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6288_ _1537_ _2901_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_88_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5088__A1 _1508_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_607 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8027_ _0236_ net1 mod.Data_Mem.F_M.MRAM\[16\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_102_255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5239_ mod.Data_Mem.F_M.MRAM\[773\]\[4\] mod.Data_Mem.F_M.MRAM\[772\]\[4\] _1903_
+ _1904_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_57_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6380__S0 _1915_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_151_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_879 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5260__A1 _1917_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_24_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_710 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_169_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_52_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_256 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__5938__I1 mod.Data_Mem.F_M.MRAM\[17\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_278 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_157_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_130_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_1061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_1094 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_153_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6512__A1 _2696_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7893__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6115__I1 mod.Data_Mem.F_M.MRAM\[6\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8249__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6019__B _2634_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_643 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8399__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_784 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_43_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5003__A1 _1552_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7565__S _3759_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4610_ _1201_ _1257_ _1281_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5590_ _1600_ _2227_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_102_1213 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4541_ _0637_ mod.Arithmetic.CN.I_in\[37\] _1213_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5085__S _1701_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6503__A1 _3106_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7260_ _3592_ _0349_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4472_ _1039_ _1144_ _1145_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__7551__I0 _3718_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6201__C _2775_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_132_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6211_ _1706_ _1794_ _2826_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_7191_ _3527_ mod.Data_Mem.F_M.MRAM\[29\]\[1\] _3550_ _3552_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_131_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6909__S _3376_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_710 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6142_ _2703_ _2757_ _2758_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_112_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7303__I0 _3618_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_765 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6708__I _3255_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6073_ mod.Data_Mem.F_M.MRAM\[797\]\[0\] _2689_ _2690_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_787 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5024_ _1579_ _1692_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_57_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1909 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6975_ _3424_ _0232_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_54_879 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7782__A3 _3446_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5926_ mod.Data_Mem.F_M.MRAM\[770\]\[4\] mod.Data_Mem.F_M.MRAM\[771\]\[4\] _2339_
+ _2547_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_41_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_710 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1087 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_146_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_55_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5857_ _2383_ mod.Data_Mem.F_M.MRAM\[773\]\[2\] _2480_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_139_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4808_ _0625_ _1367_ _1368_ _1381_ _1478_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_8576_ _0592_ net1 mod.Instr_Mem.instruction\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_166_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5788_ _1490_ _2117_ _2413_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_119_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7527_ _3744_ _3745_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_4739_ _1334_ _1343_ _1408_ _1409_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_135_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7458_ _3702_ _0437_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__7542__I0 _3754_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6409_ _2171_ mod.Data_Mem.F_M.MRAM\[12\]\[0\] _3018_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_7389_ mod.Data_Mem.F_M.MRAM\[774\]\[3\] _3668_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_122_339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_131_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_1016 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_765 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_1196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xtiny_user_project_106 la_data_out[27] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XANTENNA__4808__A1 _0625_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xtiny_user_project_117 la_data_out[38] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_29_320 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtiny_user_project_128 la_data_out[49] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_139 la_data_out[60] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_29_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8541__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5678__B _2259_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_356 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3977__I _0653_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6430__B1 _3037_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4074__S _0703_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4587__A3 _1258_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_1178 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6733__A1 mod.Data_Mem.F_M.dest\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_114_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_4_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8071__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_1127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5432__I _2086_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5311__I2 _1973_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_971 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5472__A1 _1951_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_278 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_816 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6263__I _1737_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6760_ mod.Data_Mem.F_M.MRAM\[8\]\[3\] _3287_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_62_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3972_ _0631_ _0648_ _0649_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__5775__A2 mod.Data_Mem.F_M.MRAM\[788\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5711_ _2129_ mod.Data_Mem.F_M.MRAM\[797\]\[6\] _2338_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_93_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6691_ _3242_ _3243_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6024__I0 mod.Data_Mem.F_M.MRAM\[2\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8430_ _0526_ net1 mod.Data_Mem.F_M.MRAM\[791\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5642_ _2264_ mod.Data_Mem.F_M.MRAM\[797\]\[1\] _2274_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_148_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8361_ _0457_ net1 mod.Data_Mem.F_M.MRAM\[782\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5573_ _2210_ _2211_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6212__B _2775_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7312_ _3622_ _3625_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__8414__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4524_ _1165_ _1187_ _1195_ _1196_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
X_8292_ _0388_ net1 mod.Data_Mem.F_M.MRAM\[772\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__7524__I0 _3731_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_1185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7243_ _3582_ _0342_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_102_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4455_ _0640_ mod.Arithmetic.ACTI.x\[4\] _1128_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_160_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7174_ _3542_ _0313_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4386_ _0806_ mod.Arithmetic.CN.I_in\[20\] _1059_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__4502__A3 mod.Arithmetic.CN.I_in\[20\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8564__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_540 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_713 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6125_ _2696_ _1497_ _2737_ _2741_ _1625_ _2742_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XTAP_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_584 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6056_ _2672_ _2673_ _2674_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_61_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3108 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3119 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5007_ _1514_ _1675_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_67_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2407 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2418 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_930 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_1123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2429 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1717 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1728 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_462 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_82_985 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1739 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6958_ _3397_ mod.Data_Mem.F_M.MRAM\[15\]\[3\] _3409_ _3413_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__5766__A2 _2389_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5909_ _2117_ _2531_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6889_ mod.Data_Mem.F_M.MRAM\[4\]\[4\] _3367_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_50_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5945__C _2565_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5518__A2 _2093_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_167_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_8559_ _0063_ net1 mod.Data_Mem.F_M.out_data\[23\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__5517__I _2157_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8094__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7515__I0 _3711_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_162_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_108_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_155_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_155_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtiny_user_project_12 io_oeb[1] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_1_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xtiny_user_project_23 io_oeb[12] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_77_724 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xtiny_user_project_34 io_oeb[23] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_76_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5129__S1 _1795_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xtiny_user_project_45 io_oeb[34] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XANTENNA__7931__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xtiny_user_project_56 io_out[7] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_67 io_out[26] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_78 io_out[37] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_58_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4257__A2 _0929_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xtiny_user_project_89 la_data_out[10] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_92_716 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6284__S _2044_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_429 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_91_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_610 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_40_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2930 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2941 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4009__A2 mod.Arithmetic.I_out\[73\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5206__A1 _1870_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2952 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2963 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_17_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2974 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2985 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2996 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_32_359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_158_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_38_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8437__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4193__A1 _0639_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_154_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6309__I1 _1979_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8587__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_153_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4240_ _0807_ _0915_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_99_359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5693__A1 _2321_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_101_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_68_713 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4171_ _0665_ _0842_ _0846_ _0847_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_67_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5445__A1 _2078_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7930_ _0156_ net1 mod.Data_Mem.F_M.MRAM\[8\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_49_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5996__A2 _2013_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7861_ _3917_ _3919_ _0611_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_36_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6812_ mod.Data_Mem.F_M.MRAM\[789\]\[1\] _3325_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_50_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7792_ _3888_ _3894_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__5748__A2 _1533_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6796__I1 _3312_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6743_ _3246_ mod.Data_Mem.F_M.MRAM\[0\]\[3\] _3274_ _3278_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_3955_ _0613_ _0632_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_56_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_17_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4420__A2 mod.Arithmetic.CN.I_in\[35\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_1037 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6674_ _3227_ _3228_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_149_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8413_ _0509_ net1 mod.Data_Mem.F_M.MRAM\[788\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5625_ _1845_ _2258_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__4184__A1 _0748_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8344_ _0440_ net1 mod.Data_Mem.F_M.MRAM\[780\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5556_ _1639_ _2195_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_3_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_105_615 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4507_ _0632_ _1178_ _1064_ _1070_ _1179_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_8275_ _0371_ net1 mod.Data_Mem.F_M.MRAM\[770\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5487_ _2072_ _2132_ _2133_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5273__S _1783_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7226_ _3572_ _0335_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__7954__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4438_ _1109_ _1110_ _1111_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_99_860 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_1122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7157_ _3531_ mod.Data_Mem.F_M.MRAM\[12\]\[3\] _3525_ _3532_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_115_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4369_ _0952_ _0975_ _1041_ _1042_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_59_746 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_1177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6108_ _1640_ _2722_ _2724_ _2715_ _2725_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_101_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_7088_ mod.Data_Mem.F_M.MRAM\[21\]\[7\] _3491_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_101_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6039_ _2288_ mod.Data_Mem.F_M.MRAM\[773\]\[7\] _2657_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_73_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5800__I _1612_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5987__A2 _2605_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2204 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2215 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2226 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2237 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1503 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2248 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_21 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_42_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2259 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1514 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_32 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6832__S _3337_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_43 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1536 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_54 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1547 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6787__I1 _3306_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_65 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_76 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_14_348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5295__S0 _1745_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1558 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_35_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_977 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1569 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_87 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_98 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__8090__RN net2 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_10_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6164__A2 _1702_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_163_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_135_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_123_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_819 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_151_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_607 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5675__A1 _2076_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6219__A3 mod.Data_Mem.F_M.MRAM\[20\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5427__A1 _1802_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6806__I net10 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5978__A2 mod.Data_Mem.F_M.MRAM\[782\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_546 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_643 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_1151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6490__I3 _1870_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_462 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2760 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_32_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2771 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2782 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_75_1059 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2793 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_127_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_61_977 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4402__A2 _1074_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_159_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6155__A2 _1656_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5410_ _1595_ _2069_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4166__A1 _0807_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7977__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6390_ _2252_ _2255_ _2996_ _2999_ _1489_ _2750_ _3000_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_126_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4996__I _1663_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_5341_ mod.Data_Mem.F_M.MRAM\[773\]\[6\] mod.Data_Mem.F_M.MRAM\[772\]\[6\] _1906_
+ _2004_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_138_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5093__S _1759_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8060_ _0269_ net1 mod.Data_Mem.F_M.MRAM\[20\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_114_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5272_ _1932_ mod.Data_Mem.F_M.MRAM\[789\]\[5\] _1935_ _1936_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_86_1188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4469__A2 _1141_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5666__A1 _2290_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7011_ _3227_ _3445_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_87_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5106__B _1651_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4223_ _0656_ _0831_ _0898_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_102_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_141_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4154_ _0827_ _0829_ _0830_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_56_716 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4085_ _0759_ _0760_ _0761_ _0762_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_55_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5969__A2 mod.Data_Mem.F_M.MRAM\[4\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7913_ _0139_ net1 mod.Data_Mem.F_M.MRAM\[10\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_55_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_1213 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7748__S _3867_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_7844_ _3924_ _0600_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_52_933 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_169_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7775_ _3884_ _0572_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4987_ _1584_ _1655_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__8072__RN net2 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6726_ _3266_ _0141_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_3938_ _0615_ _0616_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_6657_ mod.Data_Mem.F_M.MRAM\[27\]\[0\] _3219_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_109_217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6146__A2 _1637_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7194__I1 mod.Data_Mem.F_M.MRAM\[29\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4157__A1 _0655_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5608_ _2225_ _2240_ _2243_ _2177_ _0045_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XANTENNA__4900__S _1568_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6588_ mod.I_addr\[6\] _3183_ _3184_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__6941__I1 mod.Data_Mem.F_M.MRAM\[14\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8327_ _0423_ net1 mod.Data_Mem.F_M.MRAM\[776\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_3_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_145_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_3_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5539_ _2086_ _2179_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_105_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7282__I _3297_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8258_ _0354_ net1 mod.Data_Mem.F_M.MRAM\[5\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_106_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8132__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7209_ _3523_ mod.Data_Mem.F_M.MRAM\[2\]\[0\] _3562_ _3563_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_120_426 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8189_ _0299_ net1 mod.Data_Mem.F_M.MRAM\[19\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_115_1042 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_8_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5409__A1 _2063_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_98_1004 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5530__I _1782_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_546 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8282__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6082__A1 mod.Data_Mem.F_M.MRAM\[13\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2001 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6082__B2 mod.Data_Mem.F_M.MRAM\[12\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2012 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2023 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4632__A2 _1214_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2034 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_160_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_43_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1300 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2045 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1311 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2056 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1322 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2067 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1333 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2078 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2089 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_977 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1355 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1366 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_465 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1377 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1388 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1399 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4396__A1 _0615_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5593__B1 mod.Data_Mem.F_M.MRAM\[30\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_168_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6137__A2 mod.Data_Mem.F_M.MRAM\[14\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6932__I1 mod.Data_Mem.F_M.MRAM\[14\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4699__A2 mod.Arithmetic.CN.I_in\[69\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5896__A1 _2510_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5896__B2 _2517_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6696__I0 _3246_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6737__S _3274_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4320__A1 _0922_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_77_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_168_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_65_535 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6073__A1 mod.Data_Mem.F_M.MRAM\[797\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_80_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5820__A1 _2435_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4910_ _1578_ _1579_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_33_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5890_ _1513_ _2512_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_2590 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4841_ _1509_ _1510_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_61_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6271__I _2837_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8005__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7560_ _3766_ _0475_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4772_ mod.Arithmetic.CN.I_in\[55\] _1441_ _1442_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_140_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6511_ _2587_ mod.Data_Mem.F_M.MRAM\[13\]\[5\] _3115_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_158_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7491_ _3640_ mod.Data_Mem.F_M.MRAM\[781\]\[2\] _3720_ _3723_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_119_548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6442_ _2499_ _3050_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5887__A1 _2506_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8155__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_146_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6373_ _1655_ _2041_ _2983_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_114_220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8112_ mod.Data_Mem.F_M.out_data\[22\] net2 net1 mod.Arithmetic.CN.I_in\[22\] vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_138_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_114_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7628__A2 _3798_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5324_ mod.Data_Mem.F_M.MRAM\[5\]\[6\] mod.Data_Mem.F_M.MRAM\[4\]\[6\] _1873_ _1987_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_88_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_8043_ _0252_ net1 mod.Data_Mem.F_M.MRAM\[18\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_88_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5255_ _1906_ mod.Data_Mem.F_M.MRAM\[786\]\[4\] _1920_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__6300__A2 _2912_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4206_ _0868_ _0870_ _0880_ _0881_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XANTENNA__4311__A1 _0897_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4311__B2 mod.Arithmetic.CN.I_in\[41\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5186_ _1647_ _1851_ _1852_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_96_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_982 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4137_ _0637_ _0813_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_83_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6064__A1 _1840_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_568 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4068_ _0734_ _0742_ _0744_ _0745_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_56_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4614__A2 _1195_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7827_ _3908_ _3913_ _3914_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_52_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_169_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7277__I mod.Data_Mem.F_M.MRAM\[5\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6367__A2 _2028_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_936 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4378__A1 _0878_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7758_ _3874_ _0565_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_11_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6114__C _2708_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6709_ _3256_ mod.Data_Mem.F_M.MRAM\[28\]\[6\] _3250_ _3257_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__7316__A1 _3612_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7689_ _3838_ _0532_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6914__I1 mod.Data_Mem.F_M.MRAM\[13\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6390__I2 _2996_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_1183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_1058 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_160_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_152_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_59_362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_93_129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5802__A1 _2425_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8028__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1130 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_163_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_31_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1152 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_63_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_76_1187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1163 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1174 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1185 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1196 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_169_982 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_129_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__8178__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5030__A2 _1673_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_156_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_128_367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6905__I1 mod.Data_Mem.F_M.MRAM\[13\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5869__A1 _2124_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5869__B2 _2490_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6530__A2 mod.Data_Mem.F_M.MRAM\[12\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_48_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4541__A1 _0637_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_903 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_152_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_914 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_936 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5371__S _1890_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_958 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5040_ _1512_ _1708_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_969 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_19_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6046__A1 _2620_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_168_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6991_ _3234_ _3433_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_93_674 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7298__S _3606_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__6841__I0 _3249_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5942_ _2560_ _2561_ _2562_ _2563_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_94_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5873_ _2101_ _2495_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_90_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7612_ _3797_ _3798_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_4824_ _1492_ _1493_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_8592_ _0608_ net1 mod.Instr_Mem.instruction\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_7543_ _3755_ _0469_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_21_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4755_ mod.Arithmetic.CN.I_in\[37\] _1423_ _1213_ _1424_ _1425_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_159_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7474_ _3712_ _0443_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_162_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4686_ _0636_ _1356_ _1357_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_6425_ _3020_ _2438_ _3033_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__6521__A2 mod.Data_Mem.F_M.MRAM\[780\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6356_ mod.Data_Mem.F_M.MRAM\[13\]\[6\] _2901_ _2201_ mod.Data_Mem.F_M.MRAM\[12\]\[6\]
+ _2966_ _2967_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_89_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5307_ mod.Data_Mem.F_M.MRAM\[1\]\[5\] _1971_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5281__S _1942_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6287_ _2879_ _2885_ _2894_ _2899_ _2900_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_103_746 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_142_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_130_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8026_ _0235_ net1 mod.Data_Mem.F_M.MRAM\[16\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5238_ _1813_ _1903_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_88_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6380__S1 _2383_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4835__A2 _1503_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_1110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5169_ _1586_ _1835_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_17_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_83_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_1018 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6832__I0 _3228_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_202 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_169_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XPHY_213 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8320__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_24_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_9_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_8_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5964__B _2583_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8470__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4771__A1 _1354_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_4_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6512__A2 mod.Data_Mem.F_M.MRAM\[12\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_134_871 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_140_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6276__A1 _2846_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4287__B1 _0808_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_1180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6086__I _2702_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5204__B _1869_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_855 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6028__A1 _1670_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_674 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_90_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_90_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6750__S _3279_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_5 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_50_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5366__S _1877_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4540_ _1208_ _1211_ _1212_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_117_816 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_157_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4471_ _1042_ _1046_ _1143_ _1144_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_85_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6503__A2 mod.Data_Mem.F_M.MRAM\[769\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6210_ _2196_ _1786_ _2739_ _2825_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__4514__A1 _1185_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7190_ _3551_ _0320_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_48_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_711 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6141_ _2192_ _2689_ _2756_ _1625_ _2757_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_97_210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_711 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_722 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_48_1075 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7303__I1 mod.Data_Mem.F_M.MRAM\[768\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_755 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6072_ _2681_ _2689_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_135_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_788 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5023_ _1690_ _1691_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_85_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_749 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6019__A1 _2558_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8343__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6974_ _3386_ mod.Data_Mem.F_M.MRAM\[16\]\[0\] _3423_ _3424_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_53_335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_1160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5925_ mod.Data_Mem.F_M.MRAM\[782\]\[4\] _1901_ _2258_ _2546_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_53_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_571 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_62_891 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_167_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8493__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5856_ _2281_ mod.Data_Mem.F_M.MRAM\[772\]\[2\] _2479_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4807_ _1324_ _1475_ _1476_ _1477_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_8575_ _0079_ net1 mod.Data_Mem.F_M.out_data\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__4053__I0 _0679_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5787_ _2379_ _2393_ _2411_ _2412_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_7526_ _3407_ _3705_ _3387_ _3744_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_4738_ _1338_ _1209_ _1337_ _1408_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_163_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7457_ mod.Data_Mem.F_M.MRAM\[778\]\[5\] _3702_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_134_123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5075__I _1524_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4669_ mod.Arithmetic.CN.I_in\[46\] _1339_ _1340_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_135_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7542__I1 mod.Data_Mem.F_M.MRAM\[783\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7491__S _3720_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6408_ _2385_ _3017_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__4505__A1 _0958_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_150_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_122_307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7388_ _3667_ _0402_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_116_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_722 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6339_ _2779_ _2948_ _2949_ _2950_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_7_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6258__A1 _2870_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5305__I0 mod.Data_Mem.F_M.MRAM\[5\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xtiny_user_project_107 la_data_out[28] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_88_287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8009_ _0218_ net1 mod.Data_Mem.F_M.MRAM\[14\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xtiny_user_project_118 la_data_out[39] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_129 la_data_out[50] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_57_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5959__B _1536_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_151_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_56_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6430__A1 _2560_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6430__B2 _2388_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4992__A1 _1608_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_157_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_40_574 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4044__I0 _0680_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6733__A2 mod.Data_Mem.F_M.dest\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8501__D _0005_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4744__A1 _0622_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_126_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_85 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_153_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6497__A1 _3047_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8216__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4347__I1 _1019_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_1220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8366__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5311__I3 _1974_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_983 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_1057 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_1068 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_677 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3971_ _0639_ _0647_ _0648_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_63_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_571 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7576__S _3773_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5710_ _2071_ _2148_ _2335_ _2336_ _2337_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_62_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6690_ net5 _3242_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_31_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7221__I0 _3569_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6024__I1 mod.Data_Mem.F_M.MRAM\[3\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5641_ _2063_ _2113_ _2262_ _2273_ _0048_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_31_574 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5096__S _1565_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4735__A1 _0625_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8360_ _0456_ net1 mod.Data_Mem.F_M.MRAM\[782\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_141_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5932__B1 _2547_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5572_ _2209_ _2210_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_145_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7311_ _3624_ _0368_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_116_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4523_ _1194_ _1195_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_8291_ _0387_ net1 mod.Data_Mem.F_M.MRAM\[772\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_117_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6488__A1 _3003_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7242_ _3537_ mod.Data_Mem.F_M.MRAM\[30\]\[6\] _3579_ _3582_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_89_1197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4454_ _0915_ mod.Arithmetic.ACTI.x\[3\] _0914_ _1127_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_104_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7173_ mod.Data_Mem.F_M.MRAM\[22\]\[1\] _3542_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4385_ _0616_ _0691_ mod.Arithmetic.CN.I_in\[19\] _1058_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XTAP_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6124_ _2738_ _2740_ _2741_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XTAP_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_59_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_574 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6055_ mod.Data_Mem.F_M.MRAM\[2\]\[7\] mod.Data_Mem.F_M.MRAM\[3\]\[7\] _1769_ _2673_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_86_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_596 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5999__B1 _2611_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3109 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5006_ _1598_ _1674_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_85_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_674 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2408 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2419 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_1108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1707 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1718 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1729 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6957_ _3412_ _0226_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_109_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7883__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5908_ _2127_ _2355_ _2357_ _2527_ _2529_ _2362_ _2530_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_1
X_6888_ _3366_ _0203_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_14_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_22_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_872 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5839_ _2456_ _2462_ _2463_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_22_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_894 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__8239__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5923__B1 _2543_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4726__B2 _1273_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8558_ _0062_ net1 mod.Data_Mem.F_M.out_data\[22\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_135_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_1204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7509_ _3718_ mod.Data_Mem.F_M.MRAM\[782\]\[0\] _3734_ _3735_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_8489_ _0585_ net1 mod.Data_Mem.F_M.MRAM\[7\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_120_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5734__S _2358_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6479__A1 _3083_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_151_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_123_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8389__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtiny_user_project_13 io_oeb[2] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_24 io_oeb[13] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_49_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xtiny_user_project_35 io_oeb[24] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_77_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xtiny_user_project_46 io_oeb[35] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_118_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xtiny_user_project_57 io_out[8] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_68 io_out[27] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_76_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xtiny_user_project_79 la_data_out[0] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_76_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_45_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_942 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2920 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_84_290 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_249 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2931 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_17_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2942 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5206__A2 _1673_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6403__A1 _2422_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2953 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5201__C _1866_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2964 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2975 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4265__I0 _0768_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2986 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2997 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7203__I0 _3537_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6313__B _2873_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_127_933 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_114_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_113_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5443__I _1548_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_1023 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5693__A2 mod.Data_Mem.F_M.MRAM\[796\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4170_ _0663_ _0845_ _0846_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_122_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_1045 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_1094 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_45_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_68_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5445__A2 _2093_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_48_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7860_ _3917_ _0609_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_64_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7198__A2 _3550_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6811_ _3324_ _0168_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_51_603 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7791_ _3893_ _0579_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_35_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_63_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_51_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6742_ _3277_ _0146_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_56_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3954_ _0622_ _0630_ _0631_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_52_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6673_ net3 _3227_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_8412_ _0508_ net1 mod.Data_Mem.F_M.MRAM\[788\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5624_ _2256_ mod.Data_Mem.F_M.MRAM\[797\]\[0\] _2257_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_118_911 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_164_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8343_ _0439_ net1 mod.Data_Mem.F_M.MRAM\[778\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__8531__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5555_ _2178_ _2183_ _2194_ _0041_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_105_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4506_ mod.Arithmetic.CN.I_in\[29\] _1178_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_8274_ _0370_ net1 mod.Data_Mem.F_M.MRAM\[770\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_133_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5486_ _1799_ _2075_ _2132_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_117_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7225_ _3539_ mod.Data_Mem.F_M.MRAM\[2\]\[7\] _3567_ _3572_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_160_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4437_ _0993_ _0999_ _1110_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_28_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7156_ _3245_ _3531_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_59_714 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4368_ _0901_ _1040_ _1041_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_98_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_213 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6107_ _2723_ _1569_ _2724_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_100_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7087_ _3490_ _0278_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_63_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4299_ _0716_ _0816_ _0882_ _0709_ _0973_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_86_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_393 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_717 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6038_ mod.Data_Mem.F_M.MRAM\[770\]\[7\] mod.Data_Mem.F_M.MRAM\[771\]\[7\] _2339_
+ _2656_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_58_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2205 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_398 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2216 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2227 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2238 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6117__C _2733_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_975 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2249 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_11 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1504 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_22 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_54_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1515 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_33 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1526 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_44 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_7989_ mod.Instr_Mem.instruction\[22\] net2 net1 mod.Data_Mem.F_M.src\[0\] vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XTAP_1537 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_55 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1548 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__5295__S1 _1822_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1559 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_77 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_30_809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8061__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_168_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_148_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_88 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_41_157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_99 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_10_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_680 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5528__I _1713_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_167_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_588 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_108_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_1078 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_1201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5675__A2 _2304_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_1212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_2_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_49_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5427__A2 _2082_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_588 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_290 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3989__A2 _0665_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_569 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8404__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2750 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2761 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_166_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2772 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2783 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6822__I mod.Data_Mem.F_M.MRAM\[789\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2794 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_158_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_32_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_13_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8554__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_146_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_1082 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5340_ mod.Data_Mem.F_M.MRAM\[771\]\[6\] mod.Data_Mem.F_M.MRAM\[770\]\[6\] _1836_
+ _2003_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_115_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_1213 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_142_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6269__I _2881_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5271_ _1933_ _1934_ _1935_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_7010_ _3444_ _0247_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_114_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4222_ mod.Arithmetic.CN.I_in\[42\] _0897_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5666__A2 _2124_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4153_ _0828_ _0820_ mod.Arithmetic.CN.I_in\[33\] _0829_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_96_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4084_ _0744_ _0761_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_3_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6218__B _2508_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4517__I mod.Arithmetic.CN.I_in\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7912_ _0138_ net1 mod.Data_Mem.F_M.MRAM\[10\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__8084__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7843_ mod.Data_Mem.F_M.MRAM\[9\]\[0\] _3924_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_63_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_93_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_145_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6732__I _3234_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_1149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7774_ _3778_ mod.Data_Mem.F_M.MRAM\[797\]\[4\] _3883_ _3884_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4986_ _1638_ _1643_ _1652_ _1653_ _1654_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_51_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6725_ mod.Data_Mem.F_M.MRAM\[10\]\[5\] _3266_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_51_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3937_ _0614_ _0615_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_149_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6656_ _3218_ _0119_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__7921__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_165_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5607_ mod.Data_Mem.F_M.MRAM\[797\]\[5\] _2221_ _1749_ mod.Data_Mem.F_M.MRAM\[796\]\[5\]
+ _2242_ _2243_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XANTENNA__5354__A1 _1704_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4157__A2 mod.Arithmetic.CN.I_in\[40\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6587_ _3178_ mod.I_addr\[5\] _3179_ _3183_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_117_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8326_ _0422_ net1 mod.Data_Mem.F_M.MRAM\[776\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_30_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5538_ _2177_ _2178_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5106__A1 _1603_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8257_ _0353_ net1 mod.Data_Mem.F_M.MRAM\[5\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_65_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_755 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5469_ _2116_ _1626_ _2117_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_7208_ _3561_ _3562_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_132_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8188_ _0298_ net1 mod.Data_Mem.F_M.MRAM\[19\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__5901__I0 mod.Data_Mem.F_M.MRAM\[18\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_533 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7139_ _3508_ mod.Data_Mem.F_M.MRAM\[19\]\[5\] _3518_ _3520_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_101_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8427__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5409__A2 _0010_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_674 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6128__B _2744_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_28_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6082__A2 _2087_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2002 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2013 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_901 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2024 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2035 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1301 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2046 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8577__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2057 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1323 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2068 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1334 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2079 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1345 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_153_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1356 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1367 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1378 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1389 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5593__A1 _1953_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4396__A2 _0958_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_1093 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_155_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_6_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5896__A2 _2514_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_722 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_108_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_151_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_617 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6696__I1 mod.Data_Mem.F_M.MRAM\[28\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_1004 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_81_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4320__A2 _0660_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_801 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_717 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_78_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_77_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6073__A2 _2689_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_355 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_93_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5820__A2 _2437_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7648__I mod.Data_Mem.F_M.MRAM\[790\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_753 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4840_ _1502_ _1509_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_2580 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2591 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7944__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_1111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_159_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_33_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5584__A1 _2138_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1890 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4771_ _1354_ mod.Arithmetic.CN.I_in\[54\] _1441_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5168__I _1663_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5584__B2 _2088_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7584__S _3779_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6510_ _1966_ _3100_ _3103_ _3110_ _3114_ _0076_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai32_1
XFILLER_105_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7490_ _3722_ _0449_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_147_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4139__A2 _0814_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6441_ _2092_ _3049_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5887__A2 mod.Data_Mem.F_M.MRAM\[783\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6372_ _2882_ _2980_ _2981_ _2898_ _2078_ _2982_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_115_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8111_ mod.Data_Mem.F_M.out_data\[21\] net2 net1 mod.Arithmetic.CN.I_in\[21\] vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_5323_ mod.Data_Mem.F_M.MRAM\[15\]\[6\] _1673_ _1986_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_8042_ _0251_ net1 mod.Data_Mem.F_M.MRAM\[18\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_115_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5254_ mod.Data_Mem.F_M.MRAM\[787\]\[4\] _1919_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_87_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_69_820 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_25_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4205_ _0878_ _0879_ _0880_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_151_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4311__A2 _0833_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5631__I _1840_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5185_ mod.Data_Mem.F_M.MRAM\[770\]\[3\] _1851_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_96_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_110_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_1148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4136_ _0639_ _0811_ _0812_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_83_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_823 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6064__A2 _2402_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4247__I mod.Arithmetic.CN.I_in\[58\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_84_867 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4067_ mod.Arithmetic.CN.I_in\[15\] _0705_ _0740_ _0743_ _0744_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_84_878 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_1000 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_24_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5279__S _1942_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7558__I _3308_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_1093 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_1055 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7826_ mod.I_addr\[3\] _3911_ _3913_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_58_1066 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_169_427 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_58_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_1009 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4969_ mod.Data_Mem.F_M.MRAM\[5\]\[1\] mod.Data_Mem.F_M.MRAM\[4\]\[1\] _1636_ _1637_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_7757_ _3806_ mod.Data_Mem.F_M.MRAM\[796\]\[5\] _3872_ _3874_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_6708_ _3255_ _3256_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_22_23 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7688_ mod.Data_Mem.F_M.MRAM\[792\]\[4\] _3838_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__7316__A2 _3623_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6639_ mod.Data_Mem.F_M.MRAM\[26\]\[7\] _3210_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_20_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_106_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_1151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8309_ _0405_ net1 mod.Data_Mem.F_M.MRAM\[774\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_105_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_606 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_1195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_714 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_121_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7967__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3996__I mod.Arithmetic.ACTI.x\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1120 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1142 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1153 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1164 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7555__A2 _3762_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_85 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_1199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5566__A1 _1664_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1175 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1197 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_168_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_169_994 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_1213 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6748__S _3279_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4541__A2 mod.Arithmetic.CN.I_in\[37\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_574 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_904 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_915 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_926 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_83_1159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_948 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_959 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5451__I _1535_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7618__I0 _3749_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_823 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_569 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_878 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6990_ _3432_ _0239_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_66_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6841__I1 mod.Data_Mem.F_M.MRAM\[769\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5941_ _2256_ mod.Data_Mem.F_M.MRAM\[20\]\[4\] _2562_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_46_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_34_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6282__I _2881_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5872_ _2085_ _2484_ _2494_ _1498_ _0058_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XANTENNA__6215__C _2743_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7611_ _3296_ _3604_ _3758_ _3797_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_4823_ mod.Data_Mem.F_M.src\[1\] _1492_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_21_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8122__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8591_ _0607_ net1 mod.Data_Mem.F_M.MRAM\[9\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__5827__S _1954_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7542_ _3754_ mod.Data_Mem.F_M.MRAM\[783\]\[5\] _3752_ _3755_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4754_ _1185_ _1423_ _1424_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5309__A1 _1769_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7473_ _3711_ mod.Data_Mem.F_M.MRAM\[780\]\[3\] _3707_ _3712_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_135_806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_1015 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4685_ mod.Arithmetic.CN.I_in\[54\] _1355_ _1356_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_135_817 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5626__I _2216_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4530__I mod.Arithmetic.CN.I_in\[44\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__8272__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6424_ _2447_ _2278_ _3030_ _2420_ _2427_ _3031_ _3032_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_146_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_162_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6355_ _2903_ _2965_ _2966_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_103_703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5306_ mod.Data_Mem.F_M.MRAM\[7\]\[5\] mod.Data_Mem.F_M.MRAM\[6\]\[5\] _1515_ _1970_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_88_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6286_ _2895_ _2896_ _2897_ _2898_ _1866_ _2899_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_0_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_102_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_8025_ _0234_ net1 mod.Data_Mem.F_M.MRAM\[16\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5237_ _1901_ _1699_ _1902_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_103_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4296__A1 _0965_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7609__I0 _3784_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5168_ _1663_ _1834_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_111_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7489__S _3720_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_290 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4119_ _0672_ _0673_ _0795_ mod.P2.Rout_reg\[0\] _0796_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_84_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5099_ _1708_ _1765_ _1766_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_95_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5096__I0 _1761_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5796__A1 _2417_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7288__I _3608_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_214 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_52_561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_225 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_80_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6125__C _1625_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_7809_ mod.Data_Mem.F_M.MRAM\[7\]\[4\] _3903_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_80_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_24_285 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_71_1030 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_169_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_166_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_158_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_116_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_165_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_891 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5720__A1 _2345_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_152_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_79_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4287__A1 _0915_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_66_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_85 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_1192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6028__A2 _2118_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_62_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_165_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8145__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5787__A1 _2379_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_31_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8295__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__6051__B _2354_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4762__A2 _1429_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_117_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7000__I1 mod.Data_Mem.F_M.MRAM\[17\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4470_ _1047_ _1084_ _1142_ _1143_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_128_187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5711__A1 _2129_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4514__A2 _1093_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_131_319 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_500 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6140_ _2750_ _2755_ _2756_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_98_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_48_1087 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_745 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_609 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6071_ _2172_ _2687_ _1729_ _2688_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4278__A1 _0881_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5022_ _1522_ _1690_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_85_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_789 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_78_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6019__A2 _2631_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6424__C1 _2427_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6973_ _3422_ _3423_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_65_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1045 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6941__S _3400_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1056 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5924_ _2535_ _2140_ _2536_ _2538_ _2544_ _2545_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_59_1172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_55_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5855_ mod.Data_Mem.F_M.MRAM\[782\]\[2\] mod.Data_Mem.F_M.MRAM\[783\]\[2\] _2398_
+ _2478_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_55_1058 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4806_ _1327_ _1386_ _1476_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_8574_ _0078_ net1 mod.Data_Mem.F_M.out_data\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5786_ _2401_ _2409_ _2410_ _2411_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_148_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7525_ _3743_ _0463_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_21_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5950__A1 _2266_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4737_ _1350_ _1362_ _1407_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_107_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7456_ _3701_ _0436_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_107_327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4668_ _1203_ _1338_ _0984_ _1339_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_147_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4505__A2 _1176_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6407_ _3003_ _3008_ _3015_ _3016_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_163_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6750__I0 _3256_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5702__A1 _2203_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8018__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7387_ mod.Data_Mem.F_M.MRAM\[774\]\[2\] _3667_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__7571__I _3772_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4599_ _1152_ _1259_ _1270_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_134_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6338_ _1941_ _2002_ _2949_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_89_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_1_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_907 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5305__I1 mod.Data_Mem.F_M.MRAM\[4\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6269_ _2881_ _2882_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_48_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_8008_ _0217_ net1 mod.Data_Mem.F_M.MRAM\[14\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xtiny_user_project_108 la_data_out[29] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_119 la_data_out[40] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_57_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8168__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_951 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6415__C1 _3009_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6430__A2 _2437_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7998__RN net2 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4441__A1 _0616_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_73_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4992__A2 _1659_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5941__A1 _2256_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_5_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8175__RN net2 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6741__I0 _3243_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_69_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_79_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6097__I _2713_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4680__A1 _1227_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_169_1153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_169_1197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7989__RN net2 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3970_ _0644_ _0646_ _0647_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_63_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_391 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7221__I1 mod.Data_Mem.F_M.MRAM\[2\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5640_ _2084_ _2263_ _2272_ _2273_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XANTENNA__6185__A1 _1834_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5571_ _1548_ _2209_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_106_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5932__A1 _2423_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4735__A2 _1404_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_1110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_163_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5932__B2 _2464_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4522_ _1188_ _1193_ _1194_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_7310_ _3603_ mod.Data_Mem.F_M.MRAM\[770\]\[0\] _3623_ _3624_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_129_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8290_ _0386_ net1 mod.Data_Mem.F_M.MRAM\[772\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_89_1154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_1165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_1078 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7241_ _3581_ _0341_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__8166__RN net2 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4453_ mod.Arithmetic.CN.I_in\[65\] _1012_ _0645_ mod.Arithmetic.ACTI.x\[2\] _1126_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XFILLER_145_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_617 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4948__C _1616_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7172_ _3541_ _0312_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4384_ _1054_ _1056_ _1057_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_98_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8310__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6123_ _1795_ _1516_ _1520_ _1713_ _2739_ _2740_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XTAP_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_575 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6054_ _2495_ _2672_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_39_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5999__B2 _2613_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5005_ _1672_ _1673_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_67_951 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_569 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8460__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4671__A1 _1338_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2409 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1708 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7767__S _3878_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1719 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4255__I mod.Arithmetic.CN.I_in\[49\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_6956_ _3395_ mod.Data_Mem.F_M.MRAM\[15\]\[2\] _3409_ _3412_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_53_166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4423__A1 _0654_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5907_ mod.Data_Mem.F_M.MRAM\[16\]\[3\] mod.Data_Mem.F_M.MRAM\[17\]\[3\] _2528_ _2529_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_6887_ mod.Data_Mem.F_M.MRAM\[4\]\[3\] _3366_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_22_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5838_ _2457_ _2461_ _1804_ _2462_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_33_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_1180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_155_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5923__A1 _2539_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4726__A2 _1388_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8557_ _0061_ net1 mod.Data_Mem.F_M.out_data\[21\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_136_901 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5923__B2 _2435_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5769_ _2380_ _2394_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_7508_ _3733_ _3734_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_108_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8488_ _0584_ net1 mod.Data_Mem.F_M.MRAM\[7\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_30_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_1216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6479__A2 _1855_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8157__RN net2 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_146_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7439_ mod.Data_Mem.F_M.MRAM\[777\]\[4\] _3693_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__7007__S _3440_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_77_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xtiny_user_project_14 io_oeb[3] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_77_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xtiny_user_project_25 io_oeb[14] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_36 io_oeb[25] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_49_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtiny_user_project_47 io_oeb[36] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_77_748 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xtiny_user_project_58 io_out[9] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_103_396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xtiny_user_project_69 io_out[28] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_40_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_92_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_461 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4662__A1 mod.Arithmetic.CN.I_in\[38\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2910 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2921 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2932 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_75_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2943 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7600__A1 _1787_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6403__A2 _3010_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2954 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2965 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4414__A1 _0992_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2976 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4265__I1 _0773_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4414__B2 _0988_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2987 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_32_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2998 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_13_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7203__I1 mod.Data_Mem.F_M.MRAM\[29\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6167__A1 _2708_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_145_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5925__S _2258_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_127_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__8333__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8148__RN net2 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_45_1057 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8483__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4653__A1 _1285_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7587__S _3779_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_965 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4075__I _0630_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6810_ mod.Data_Mem.F_M.MRAM\[789\]\[0\] _3324_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_35_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_24_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_63_464 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4405__A1 _0620_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7790_ _3309_ mod.Data_Mem.F_M.MRAM\[798\]\[3\] _3889_ _3893_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__5602__B1 mod.Data_Mem.F_M.MRAM\[30\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6741_ _3243_ mod.Data_Mem.F_M.MRAM\[0\]\[2\] _3274_ _3277_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_50_125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3953_ mod.Arithmetic.CN.I_in\[8\] _0630_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6504__B _2474_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_1153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6290__I _1564_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_52_1017 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6672_ _3226_ _0127_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_31_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8411_ _0507_ net1 mod.Data_Mem.F_M.MRAM\[788\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5623_ _2060_ _2256_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5835__S _2452_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8342_ _0438_ net1 mod.Data_Mem.F_M.MRAM\[778\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5554_ _2184_ _2193_ _2194_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4505_ _0958_ _1176_ _1177_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__8139__RN net2 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6705__I0 _3253_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5485_ _2129_ mod.Data_Mem.F_M.MRAM\[799\]\[3\] _2130_ _2131_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_8273_ _0369_ net1 mod.Data_Mem.F_M.MRAM\[770\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_105_617 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5634__I _1493_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7224_ _3571_ _0334_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4436_ _0930_ _0995_ _0996_ _0997_ _0994_ _1109_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_99_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_7155_ _3530_ _0306_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4367_ _0970_ _0974_ _1040_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_86_501 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4892__A1 _1554_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_1157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6106_ _1737_ _2723_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_7086_ mod.Data_Mem.F_M.MRAM\[21\]\[6\] _3490_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_58_225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7130__I0 _3450_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4298_ _0971_ _0972_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__4694__B _1364_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_383 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_394 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6094__B1 mod.Data_Mem.F_M.MRAM\[791\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_355 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6037_ mod.Data_Mem.F_M.MRAM\[782\]\[7\] mod.Data_Mem.F_M.MRAM\[783\]\[7\] _2326_
+ _2655_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_100_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4644__A1 _1063_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2206 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2217 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2228 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7497__S _3726_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2239 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_12 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_55_987 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1505 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8206__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_23 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1516 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_7988_ mod.Instr_Mem.instruction\[17\] net2 net1 mod.P1.instr_reg\[17\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XTAP_1527 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_45 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1538 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_56 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_42_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_1220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_67 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1549 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6939_ _3399_ mod.Data_Mem.F_M.MRAM\[14\]\[4\] _3400_ _3401_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XPHY_78 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_23_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_161_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6133__C _2084_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8356__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_168_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6944__I0 _3403_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4580__B1 _1136_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5544__I _1804_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_151_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_123_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_2_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4183__I0 _0748_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_49_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_85 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_45_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_46_987 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2740 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2751 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2762 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2773 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2784 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2795 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5719__I _1714_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5060__A1 _1631_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_1050 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_398 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6560__A1 _2831_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_753 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_51_1094 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5270_ mod.Data_Mem.F_M.MRAM\[788\]\[5\] _1934_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__6312__A1 _2870_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7873__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4221_ _0643_ mod.Arithmetic.CN.I_in\[42\] _0896_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_68_501 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_832 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4152_ _0618_ _0828_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__7112__I0 _3452_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6285__I _2837_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4083_ _0736_ _0741_ _0760_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__8229__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4626__A1 _1293_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7911_ _0137_ net1 mod.Data_Mem.F_M.MRAM\[10\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_48_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7842_ _3923_ _0599_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6379__A1 _2886_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7110__S _3501_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8379__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7773_ _3877_ _3883_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_168_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_52_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5051__A1 _1713_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4985_ _1556_ _1653_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6724_ _3265_ _0140_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_3936_ _0613_ _0614_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_32_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6926__I0 _3386_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6655_ mod.Data_Mem.F_M.MRAM\[25\]\[7\] _3218_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_164_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5606_ _1940_ _2241_ _2242_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__5354__A2 _2016_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6551__A1 _2511_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4157__A3 mod.Arithmetic.CN.I_in\[41\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6586_ _3182_ _0085_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_118_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8325_ _0421_ net1 mod.Data_Mem.F_M.MRAM\[776\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5537_ _2158_ _2132_ _2177_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_117_252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_105_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7780__S _3883_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8256_ _0352_ net1 mod.Data_Mem.F_M.MRAM\[5\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__6303__A1 _2870_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5106__A2 _1772_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_160_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5468_ _1812_ _2116_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_7207_ _3270_ _3272_ _3389_ _3561_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_4419_ _0893_ _0980_ _1092_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_8187_ _0297_ net1 mod.Data_Mem.F_M.MRAM\[19\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__5901__I1 mod.Data_Mem.F_M.MRAM\[19\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_99_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5399_ _2059_ _2060_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_87_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7138_ _3519_ _0300_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_101_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7069_ _3481_ _0269_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_98_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2003 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2014 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2025 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2036 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1302 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2047 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1313 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_710 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2058 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1324 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2069 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1335 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1346 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1357 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5539__I _2086_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5042__A1 _1708_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1368 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_146_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_70_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5593__A2 mod.Data_Mem.F_M.MRAM\[31\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4396__A3 _1063_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_167_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_161_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_1015 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_35_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_11_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7754__I _3866_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6542__A1 _3083_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7590__I0 _3784_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7896__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_797 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_285 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7342__I0 _3615_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_1021 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_1190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_1016 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__4320__A3 _0840_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_526 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8521__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3260 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2570 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2581 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2592 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_765 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6230__B1 _2835_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_1161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_1123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1880 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4770_ _0624_ _1439_ _1440_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_1891 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_105_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7664__I mod.Data_Mem.F_M.MRAM\[791\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_146_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_1208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6440_ _3030_ _2451_ _3046_ _2672_ _3047_ _3048_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XANTENNA__6533__A1 _2522_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5336__A2 _1998_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_162_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_61_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6371_ _2034_ _2035_ _2180_ _2981_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_115_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8110_ mod.Data_Mem.F_M.out_data\[20\] net2 net1 mod.Arithmetic.CN.I_in\[20\] vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_5322_ _1899_ _1963_ _1985_ _0005_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_142_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_103_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8041_ _0250_ net1 mod.Data_Mem.F_M.MRAM\[18\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5253_ _1779_ _1918_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_69_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8051__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4204_ _0876_ _0872_ _0874_ _0879_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
X_5184_ _1614_ _1843_ _1849_ _1850_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_69_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4135_ _0644_ _0805_ _0810_ _0811_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XANTENNA__6944__S _3400_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_898 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4066_ _0737_ _0743_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__7839__I _3169_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5272__A1 _1932_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_1083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7013__A2 _3446_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7825_ _3907_ _3912_ _0594_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_52_787 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7756_ _3873_ _0564_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_51_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_1212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4968_ _1594_ _1636_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_51_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_149_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6707_ net9 _3255_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_138_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7687_ _3837_ _0531_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4899_ _1567_ _1568_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_165_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6638_ _3209_ _0110_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6524__A1 _2500_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7572__I0 _3771_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6569_ _0612_ _3169_ _3170_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_106_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_8308_ _0404_ net1 mod.Data_Mem.F_M.MRAM\[774\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_69_1163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7324__I0 _3618_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_161_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_154_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8239_ _0335_ net1 mod.Data_Mem.F_M.MRAM\[2\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_156_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7015__S _3448_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8544__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_995 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5978__B _2597_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_27_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1110 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_1213 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1121 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1132 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_63_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5015__A1 _1681_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5269__I _1692_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1143 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1154 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1165 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1187 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1198 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_8_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7484__I _3292_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6515__A1 _3060_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7563__I0 _3754_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6515__B2 _3020_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_155_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_144_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_109_572 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8074__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_1165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_151_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_83_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_916 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_949 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_927 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_938 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_759 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_949 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7618__I1 mod.Data_Mem.F_M.MRAM\[787\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7911__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_18_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_5940_ _2326_ mod.Data_Mem.F_M.MRAM\[21\]\[4\] _2561_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_81_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3090 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5871_ _2489_ _2493_ _2494_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_34_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_61_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5179__I _1578_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7610_ _3796_ _0495_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4822_ _1490_ _1491_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_8590_ _0606_ net1 mod.Data_Mem.F_M.MRAM\[9\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_33_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7541_ _3315_ _3754_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4753_ mod.Arithmetic.CN.I_in\[38\] _1423_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_30_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6512__B _2596_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8417__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5309__A2 _1971_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7472_ _3308_ _3711_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_88_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4684_ mod.Arithmetic.CN.I_in\[52\] _1354_ _1355_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_6423_ _2388_ _3031_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6939__S _3400_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_6354_ _2134_ mod.Data_Mem.F_M.MRAM\[15\]\[6\] mod.Data_Mem.F_M.MRAM\[14\]\[6\] _2216_
+ _2965_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__7306__I0 _3620_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8567__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5305_ mod.Data_Mem.F_M.MRAM\[5\]\[5\] mod.Data_Mem.F_M.MRAM\[4\]\[5\] _1968_ _1969_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_103_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6285_ _2837_ _2898_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_88_426 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8024_ _0233_ net1 mod.Data_Mem.F_M.MRAM\[16\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5236_ mod.Data_Mem.F_M.MRAM\[783\]\[4\] _1901_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_102_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_971 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7609__I1 mod.Data_Mem.F_M.MRAM\[786\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_29_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5167_ _1764_ _1832_ _1531_ _1833_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_96_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_57_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_846 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4118_ _0794_ _0795_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_5098_ mod.Data_Mem.F_M.MRAM\[770\]\[2\] _1765_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__7569__I _3292_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5096__I1 _1762_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4049_ _0691_ _0726_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_71_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6406__C _3014_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__5089__I _1499_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6045__I0 mod.Data_Mem.F_M.MRAM\[16\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_7808_ _3902_ _0587_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XPHY_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_713 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_237 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_724 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_169_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_248 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__7793__I0 _3312_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7739_ _3863_ _0557_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_71_1053 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_162_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__8097__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6141__C _1625_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_126_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5720__A2 mod.Data_Mem.F_M.MRAM\[28\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_165_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7934__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5484__A1 _1879_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_781 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_816 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6284__I0 _1921_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5787__A2 _2393_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_646 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_70_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7784__I0 _3293_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_31_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_15_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7536__I0 _3711_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_8_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3970__A1 _0644_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_391 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5711__A2 mod.Data_Mem.F_M.MRAM\[797\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_713 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_724 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7464__A2 _3705_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6070_ _2686_ _2687_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_746 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_48_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_1058 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_757 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_718 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_24_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_5021_ _1685_ mod.Data_Mem.F_M.MRAM\[789\]\[1\] _1688_ _1689_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_79_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6424__B1 _3030_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6424__C2 _3031_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6972_ _3269_ _3270_ _3421_ _3422_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_19_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5923_ _2539_ _2541_ _2543_ _2435_ _2544_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_53_359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_540 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_1184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5854_ _2475_ _1765_ _2476_ _2477_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_21_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_107_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4805_ _1327_ _1386_ _1475_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_8573_ _0077_ net1 mod.Data_Mem.F_M.out_data\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__5637__I _1811_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5785_ _2377_ _2410_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6242__B _2738_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7524_ _3731_ mod.Data_Mem.F_M.MRAM\[782\]\[7\] _3739_ _3743_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4736_ _1293_ _1402_ _1405_ _1406_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_119_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5950__A2 mod.Data_Mem.F_M.MRAM\[4\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7455_ mod.Data_Mem.F_M.MRAM\[778\]\[4\] _3701_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_107_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4667_ mod.Arithmetic.CN.I_in\[45\] _1338_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__7957__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6406_ _2110_ _2387_ _3013_ _3014_ _3015_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_162_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7386_ _3666_ _0401_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6750__I1 mod.Data_Mem.F_M.MRAM\[0\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4598_ _1260_ _1261_ _1269_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_89_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6337_ _1635_ _2003_ _2948_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_103_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_746 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_66_1188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6268_ _2707_ _2691_ _2881_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_103_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_8007_ _0216_ net1 mod.Data_Mem.F_M.MRAM\[14\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_9_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5219_ _1653_ _1884_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xtiny_user_project_109 la_data_out[30] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_69_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6199_ _2425_ mod.Data_Mem.F_M.MRAM\[22\]\[2\] mod.Data_Mem.F_M.MRAM\[23\]\[2\] _2448_
+ _2814_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_97_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6415__B1 _3022_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_816 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6415__C2 _2368_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_646 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_1104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4441__A2 mod.Arithmetic.CN.I_in\[51\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6931__I _3242_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_166_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7518__I0 _3725_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_165_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_154_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_1200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6741__I1 mod.Data_Mem.F_M.MRAM\[0\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_85 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8112__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7203__S _3553_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__4680__A2 _1230_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7002__I _3434_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8262__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_1204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7757__I0 _3806_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_690 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5457__I _1495_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5570_ _2178_ _2199_ _2208_ _0042_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__7509__I0 _3718_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6980__I1 mod.Data_Mem.F_M.MRAM\[16\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_156_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4521_ _1190_ _1079_ _1191_ _1192_ _1193_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
X_7240_ _3569_ mod.Data_Mem.F_M.MRAM\[30\]\[5\] _3579_ _3581_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_89_1177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4452_ _0614_ mod.Arithmetic.CN.I_in\[68\] _1125_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_144_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4499__A2 _1064_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6288__I _1537_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7171_ mod.Data_Mem.F_M.MRAM\[22\]\[0\] _3541_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4383_ _0634_ _0959_ _0809_ _1055_ _1056_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XFILLER_131_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6122_ _2706_ _2739_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_113_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_112_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_532 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_716 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6053_ _2185_ _2154_ _2670_ _2263_ _2671_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_85_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_100_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_576 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5999__A2 _2150_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5004_ _1598_ _1672_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_100_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4671__A2 _1209_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_148_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_66_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1709 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6955_ _3411_ _0225_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_54_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5620__A1 _1940_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4423__A2 mod.Arithmetic.CN.I_in\[44\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5906_ _1894_ _2528_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_6886_ _3365_ _0202_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__7748__I0 _3747_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5837_ _2458_ _2454_ _2367_ _2459_ _2460_ _2170_ _2461_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XANTENNA__5908__C1 _2529_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4187__A1 _0802_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_148_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8556_ _0060_ net1 mod.Data_Mem.F_M.out_data\[20\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__5923__A2 _2541_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_1192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5768_ _2382_ _2384_ _2392_ _2393_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_120_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_7507_ _3634_ _3387_ _3389_ _3733_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_108_615 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4719_ _1273_ _1389_ _1390_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_8487_ _0583_ net1 mod.Data_Mem.F_M.MRAM\[798\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5699_ _2326_ mod.Data_Mem.F_M.MRAM\[28\]\[5\] _2259_ _2327_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_147_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7438_ _3692_ _0427_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_163_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_607 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5231__S0 _1751_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8135__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_155_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7369_ mod.Data_Mem.F_M.MRAM\[773\]\[1\] _3658_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_1_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_103_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xtiny_user_project_15 io_oeb[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_26 io_oeb[15] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_130_150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtiny_user_project_37 io_oeb[26] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_162_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xtiny_user_project_48 io_oeb[37] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XANTENNA__5830__I _2354_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8285__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6100__A2 _2689_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xtiny_user_project_59 io_out[10] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_130_183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4111__A1 _0740_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_985 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5051__B _1651_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2900 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2911 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_17_326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2922 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2933 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2944 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_17_359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2955 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2966 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5478__S _1890_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8093__RN net2 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2977 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_32_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5611__A1 mod.Data_Mem.F_M.MRAM\[29\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5611__B2 mod.Data_Mem.F_M.MRAM\[28\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2988 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2999 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_690 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5277__I _1940_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5678__A1 _2295_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_153_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_45_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_122_651 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6836__I _3336_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4102__A1 _0727_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_248 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_879 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_67_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_985 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_730 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_977 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_988 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5602__A1 _1953_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6571__I mod.I_addr\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8008__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6740_ _3276_ _0145_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_3952_ _0628_ _0629_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_95_1181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA_output8_I net8 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_1023 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6671_ mod.Data_Mem.F_M.MRAM\[27\]\[7\] _3226_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_143_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_91_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4091__I mod.Arithmetic.ACTI.x\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4169__A1 _0844_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8410_ _0506_ net1 mod.Data_Mem.F_M.MRAM\[788\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5622_ _2225_ _2252_ _2255_ _2177_ _0047_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XANTENNA__8158__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8341_ _0437_ net1 mod.Data_Mem.F_M.MRAM\[778\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_157_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5553_ _2169_ _2185_ _2159_ _2192_ _2193_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XANTENNA__7108__S _3501_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5915__I _2440_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_968 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6012__S _2418_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4504_ _0806_ _1062_ mod.Arithmetic.CN.I_in\[29\] _1176_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_8272_ _0368_ net1 mod.Data_Mem.F_M.MRAM\[770\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5484_ _1879_ mod.Data_Mem.F_M.MRAM\[798\]\[3\] _2130_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_145_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6705__I1 mod.Data_Mem.F_M.MRAM\[28\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5669__A1 _2074_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7223_ _3537_ mod.Data_Mem.F_M.MRAM\[2\]\[6\] _3567_ _3571_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__6947__S _3400_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4435_ _1000_ _1001_ _1106_ _1107_ _1004_ _1108_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai32_2
XFILLER_99_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7154_ _3529_ mod.Data_Mem.F_M.MRAM\[12\]\[2\] _3525_ _3530_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4366_ _0951_ _1037_ _1038_ _1039_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__4975__B _1642_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_59_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4892__A2 _1504_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6105_ _2620_ mod.Data_Mem.F_M.MRAM\[774\]\[0\] mod.Data_Mem.F_M.MRAM\[775\]\[0\]
+ _2162_ _2722_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_141_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_362 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_63_1169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7085_ _3489_ _0277_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4297_ _0618_ mod.Arithmetic.CN.I_in\[11\] _0971_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_112_183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6094__A1 _2326_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6094__B2 _2116_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6036_ _2535_ _2156_ _2536_ _2649_ _2653_ _2654_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_67_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7778__S _3883_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_55_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2207 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2218 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2229 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_148_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_13 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_54_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1506 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_7987_ mod.Instr_Mem.instruction\[13\] net2 net1 mod.P1.instr_reg\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XPHY_24 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_42_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1517 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_35 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__8075__RN net2 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_46 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_14_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1539 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_57 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_6938_ _3390_ _3400_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XPHY_68 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_81_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_79 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_161_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6869_ mod.Data_Mem.F_M.MRAM\[6\]\[2\] _3357_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5097__I _1607_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6944__I1 mod.Data_Mem.F_M.MRAM\[14\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_568 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8539_ _0043_ net1 mod.Data_Mem.F_M.out_data\[35\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__5825__I _2448_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7018__S _3448_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_159_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4580__A1 _1251_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4580__B2 _1017_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4332__A1 _0665_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_104_651 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_77_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5832__A1 _2447_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_538 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_793 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_432 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_166_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_57_292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2730 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2741 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2752 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2763 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2774 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2785 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2796 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8300__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_682 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6935__I1 mod.Data_Mem.F_M.MRAM\[14\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_158_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_51_1062 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5735__I _1677_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4571__A1 mod.Arithmetic.CN.I_in\[67\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8450__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_1158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6312__A2 _1950_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4220_ _0892_ _0893_ _0894_ _0895_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__4323__A1 _0653_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_971 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_123_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4151_ _0652_ _0826_ _0827_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_95_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7112__I1 mod.Data_Mem.F_M.MRAM\[3\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6076__A1 mod.Data_Mem.F_M.MRAM\[781\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_568 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4082_ _0757_ _0758_ _0732_ _0759_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_110_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_1180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7910_ _0136_ net1 mod.Data_Mem.F_M.MRAM\[10\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_97_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_730 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_64_752 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7841_ _0610_ _3922_ _3923_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_24_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7772_ _3882_ _0571_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5587__B1 _2224_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4984_ _1645_ _1648_ _1650_ _1651_ _1652_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_23_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6723_ mod.Data_Mem.F_M.MRAM\[10\]\[4\] _3265_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_3935_ mod.Arithmetic.CN.F_in\[0\] _0613_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_20_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6654_ _3217_ _0118_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6926__I1 mod.Data_Mem.F_M.MRAM\[14\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5605_ _2233_ mod.Data_Mem.F_M.MRAM\[799\]\[5\] mod.Data_Mem.F_M.MRAM\[798\]\[5\]
+ _2234_ _2241_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_118_710 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6585_ mod.I_addr\[5\] _3181_ _3182_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__6551__A2 mod.Data_Mem.F_M.MRAM\[0\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8324_ _0420_ net1 mod.Data_Mem.F_M.MRAM\[776\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_118_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_106_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5536_ _2176_ _0040_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_3_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8255_ _0351_ net1 mod.Data_Mem.F_M.MRAM\[31\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_117_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5467_ _2095_ _2099_ _2105_ _2115_ _0032_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__7860__I _3917_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7206_ _3560_ _0327_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_133_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5362__I0 mod.Data_Mem.F_M.MRAM\[1\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4418_ _0655_ _1090_ _1091_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_8186_ _0296_ net1 mod.Data_Mem.F_M.MRAM\[19\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_114_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5398_ _1522_ _2059_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_120_429 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_160_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7137_ _3456_ mod.Data_Mem.F_M.MRAM\[19\]\[4\] _3518_ _3519_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_101_610 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4349_ _0992_ _1002_ _1022_ _1023_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_86_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6067__A1 _2682_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_47_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7068_ mod.Data_Mem.F_M.MRAM\[20\]\[5\] _3481_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_74_505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4078__B1 _0708_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6019_ _2558_ _2631_ _2634_ _2637_ _2638_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_74_538 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_27_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_730 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2004 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_752 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2015 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2026 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8323__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2037 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1303 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2048 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1314 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2059 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1325 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1336 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_969 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1347 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_755 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1358 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1369 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_168_33 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_10_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__8473__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_168_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_128_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6542__A2 mod.Data_Mem.F_M.MRAM\[768\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_164_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7342__I1 mod.Data_Mem.F_M.MRAM\[771\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5290__I _1953_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6058__A1 _2062_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_974 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_80 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7211__S _3562_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3250 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3261 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_80_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_2560 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2571 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2582 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6230__A1 _2831_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2593 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6230__B2 _2093_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1870 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1881 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_980 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1892 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4792__A1 _0696_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7030__I0 _3416_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6533__A2 mod.Data_Mem.F_M.MRAM\[0\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4544__A1 _1214_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6370_ _2032_ _2033_ _1738_ _2980_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_127_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5321_ _1966_ _1984_ _1985_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_114_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6297__A1 _2752_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8040_ _0249_ net1 mod.Data_Mem.F_M.MRAM\[18\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_115_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7990__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5252_ _1700_ _1916_ _1917_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_64_1220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4203_ _0877_ _0878_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_68_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5183_ _1844_ _1848_ _1849_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_151_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6049__A1 _1612_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4134_ _0646_ _0809_ _0810_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_84_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8346__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_83_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_538 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4065_ _0736_ _0741_ _0742_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_37_752 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_83_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7549__A1 _3232_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_571 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7824_ _3907_ _3911_ _3912_ _0593_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_51_210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_1046 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8496__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_40_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7755_ _3778_ mod.Data_Mem.F_M.MRAM\[796\]\[4\] _3872_ _3873_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_52_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4967_ _1584_ _1635_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_6706_ _3254_ _0133_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4783__A1 _0743_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7686_ mod.Data_Mem.F_M.MRAM\[792\]\[3\] _3837_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4898_ _1513_ _1567_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__7021__I0 _3452_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_164_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6637_ mod.Data_Mem.F_M.MRAM\[26\]\[6\] _3209_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__8202__RN net2 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6524__A2 _2602_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6568_ mod.I_addr\[1\] _3169_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_4_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_152_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8307_ _0403_ net1 mod.Data_Mem.F_M.MRAM\[774\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5519_ _1527_ _2160_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_105_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6499_ mod.Data_Mem.F_M.MRAM\[780\]\[4\] mod.Data_Mem.F_M.MRAM\[782\]\[4\] mod.Data_Mem.F_M.MRAM\[781\]\[4\]
+ _1901_ _2270_ _3083_ _3104_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__7324__I1 mod.Data_Mem.F_M.MRAM\[770\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_1175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_1017 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8238_ _0334_ net1 mod.Data_Mem.F_M.MRAM\[2\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5335__I0 _1994_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4299__B1 _0882_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_278 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8169_ mod.Data_Mem.F_M.out_data\[79\] net2 net1 mod.Arithmetic.I_out\[79\] vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_59_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6934__I _3245_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_730 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6460__A1 _3021_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6460__B2 _3031_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_1113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_722 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_1100 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8073__D mod.P3.Res\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_21 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_1111 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1122 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1133 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1144 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6212__A1 _1734_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1155 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_163_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4074__I0 mod.Arithmetic.CN.I_in\[17\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_169_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7863__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1177 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1188 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1199 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_169_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6515__A2 _2591_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8219__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6279__A1 _2891_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_1117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5326__I0 mod.Data_Mem.F_M.MRAM\[1\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_906 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_917 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8369__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_939 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_78_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6451__A1 _2258_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3080 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3091 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5870_ _2457_ _2492_ _1804_ _2493_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_34_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4821_ _1489_ _1490_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_2390 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_574 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_7540_ _3753_ _0468_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_21_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4752_ _0623_ _1422_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_105_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7003__I0 _3399_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_146_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7471_ _3710_ _0442_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_105_1055 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4683_ mod.Arithmetic.CN.I_in\[53\] _1354_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_6422_ _2429_ _3030_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_162_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_88_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6353_ _2951_ _2954_ _2960_ _2963_ _2964_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__5190__A1 _1658_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_161_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7306__I1 mod.Data_Mem.F_M.MRAM\[768\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5304_ _1509_ _1968_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__5317__I0 mod.Data_Mem.F_M.MRAM\[17\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6284_ _1921_ _1922_ _2044_ _2897_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8023_ _0232_ net1 mod.Data_Mem.F_M.MRAM\[16\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__5868__I1 mod.Data_Mem.F_M.MRAM\[17\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5235_ _1871_ _1885_ _1887_ _1897_ _1899_ _1900_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_64_1050 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_546 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_69_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5166_ mod.Data_Mem.F_M.MRAM\[791\]\[3\] mod.Data_Mem.F_M.MRAM\[790\]\[3\] _1581_
+ _1832_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_97_983 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_151_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4117_ _0673_ _0676_ _0791_ _0793_ _0794_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_110_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5097_ _1607_ _1764_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_84_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4048_ _0724_ _0725_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_84_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7886__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7786__S _3889_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_65_891 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_24_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7242__I0 _3537_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6045__I1 mod.Data_Mem.F_M.MRAM\[17\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_216 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_24_254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_7807_ mod.Data_Mem.F_M.MRAM\[7\]\[3\] _3902_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_24_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_52_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5999_ _2535_ _2150_ _2611_ _2613_ _2617_ _2618_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XPHY_249 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__7793__I1 mod.Data_Mem.F_M.MRAM\[798\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_1021 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4756__A1 mod.Arithmetic.CN.I_in\[39\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7738_ mod.Data_Mem.F_M.MRAM\[795\]\[5\] _3863_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_71_1032 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5319__B _1508_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_165_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7669_ _3828_ _0522_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_125_307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5181__A1 _1647_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8511__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5833__I _2366_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5054__B _1721_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6130__B1 _1809_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6808__I0 mod.Data_Mem.F_M.MRAM\[799\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6028__A4 _2646_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6433__A1 _2626_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6284__I1 _1922_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_167_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7233__I0 _3529_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_714 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4912__I _1580_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8041__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_157_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7536__I1 mod.Data_Mem.F_M.MRAM\[783\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_102_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3970__A2 _0646_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8191__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5172__A1 _1834_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_1023 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_703 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_714 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_48_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_568 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5020_ _1686_ _1687_ _1688_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5475__A2 _2122_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6424__A1 _2447_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6424__B2 _2420_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6971_ _3420_ _3421_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_54_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1014 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_1130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_72 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5922_ _2151_ _1919_ _2542_ _2543_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__4986__A1 _1638_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_1152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5853_ _2161_ mod.Data_Mem.F_M.MRAM\[771\]\[2\] _2476_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__6523__B _2406_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_1106 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5918__I _2402_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_146_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_1049 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4822__I _1490_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6283__S0 _2448_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4738__A1 _1338_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4804_ _1406_ _1432_ _1473_ _1474_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
X_8572_ _0076_ net1 mod.Data_Mem.F_M.out_data\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5784_ _2405_ _2408_ _2409_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_9_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_147_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7523_ _3742_ _0462_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_21_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4735_ _0625_ _1404_ _1405_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__8534__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7454_ _3700_ _0435_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_163_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4666_ _1251_ _1336_ _1337_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_31_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6405_ _2100_ _3014_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_7385_ mod.Data_Mem.F_M.MRAM\[774\]\[1\] _3666_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4597_ mod.Arithmetic.ACTI.x\[6\] _1267_ _0796_ _1268_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_116_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6336_ _2846_ _2945_ _2946_ _2947_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_66_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_1213 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_1009 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6267_ _1889_ _1891_ _2723_ _2880_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_88_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5466__A2 _2112_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8006_ _0215_ net1 mod.Data_Mem.F_M.MRAM\[13\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5218_ _1874_ _1876_ _1878_ _1880_ _1881_ _1882_ _1883_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_57_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6198_ _2765_ _2811_ _2812_ _2813_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_130_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8525__181 net181 vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
X_5149_ mod.Data_Mem.F_M.MRAM\[3\]\[3\] mod.Data_Mem.F_M.MRAM\[1\]\[3\] mod.Data_Mem.F_M.MRAM\[0\]\[3\]
+ mod.Data_Mem.F_M.MRAM\[2\]\[3\] _1812_ _1814_ _1815_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_45_806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6415__A1 _3021_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6415__B2 _3023_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_677 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_84_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8064__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7215__I0 _3531_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5828__I _1519_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7518__I1 mod.Data_Mem.F_M.MRAM\[782\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5764__S _1581_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_20_290 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7901__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5563__I _2201_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_1212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4901__A1 _1566_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_1109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_739 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6394__I _1724_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8407__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6406__A1 _2110_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_169_1122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_169_1133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_48_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_1049 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8557__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_680 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7757__I1 mod.Data_Mem.F_M.MRAM\[796\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_533 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_393 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4520_ mod.Arithmetic.CN.I_in\[11\] _1078_ _1192_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_145_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_117_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4451_ _1008_ _1014_ _1123_ _1124_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_7_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7170_ _3540_ _0311_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4382_ _0844_ mod.Arithmetic.CN.I_in\[26\] _1055_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XTAP_500 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4089__I _0746_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6121_ _2373_ _2691_ _2738_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_112_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_533 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_544 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6052_ _2539_ _2663_ _2666_ _2669_ _2670_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XTAP_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_588 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5003_ _1552_ _1634_ _1668_ _1670_ _1671_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_152_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_61_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8087__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_677 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_38_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_1127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4959__A1 _1539_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6954_ _3393_ mod.Data_Mem.F_M.MRAM\[15\]\[1\] _3409_ _3411_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_42_809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5905_ mod.Data_Mem.F_M.MRAM\[14\]\[3\] mod.Data_Mem.F_M.MRAM\[15\]\[3\] _2331_ _2527_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_81_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6885_ mod.Data_Mem.F_M.MRAM\[4\]\[2\] _3365_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5648__I _2088_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5836_ mod.Data_Mem.F_M.MRAM\[16\]\[1\] mod.Data_Mem.F_M.MRAM\[17\]\[1\] _2152_ _2460_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_14_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7924__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4187__A2 _0818_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5767_ _2210_ _2387_ _2391_ _2392_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_8555_ _0059_ net1 mod.Data_Mem.F_M.out_data\[19\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_136_903 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7506_ _3732_ _0455_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4718_ _1276_ _1388_ _1389_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_8486_ _0582_ net1 mod.Data_Mem.F_M.MRAM\[798\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5698_ _1517_ _2326_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_68_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7437_ mod.Data_Mem.F_M.MRAM\[777\]\[3\] _3692_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_107_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4649_ _1303_ _1319_ _1320_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_162_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5231__S1 _1882_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7368_ _3657_ _0392_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_118_1021 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6319_ _1603_ _1937_ _2931_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_131_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_855 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7299_ _3616_ _0364_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xtiny_user_project_16 io_oeb[5] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_103_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtiny_user_project_27 io_oeb[16] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_77_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_588 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xtiny_user_project_38 io_oeb[27] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_49 io_out[0] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_131_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_131_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_430 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_975 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2901 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2912 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5759__S _2383_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2923 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_17_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2934 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2945 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_169_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4890__C _1551_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2956 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2967 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5611__A2 _2086_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2978 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2989 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_52_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_158_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4178__A2 _0673_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_127_936 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5127__A1 _1791_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_154_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6324__B1 mod.Data_Mem.F_M.MRAM\[14\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_1080 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_1015 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_964 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_48_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7052__A1 _3316_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_63_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7947__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5602__A2 mod.Data_Mem.F_M.MRAM\[31\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3951_ _0627_ _0628_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_50_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_44_680 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_1133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5468__I _1812_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6670_ _3225_ _0126_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_32_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5621_ mod.Data_Mem.F_M.MRAM\[797\]\[7\] _2226_ _2227_ mod.Data_Mem.F_M.MRAM\[796\]\[7\]
+ _2254_ _2255_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XFILLER_91_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4169__A2 mod.Arithmetic.ACTI.x\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_31_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6563__B1 _3107_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8340_ _0436_ net1 mod.Data_Mem.F_M.MRAM\[778\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5552_ mod.Data_Mem.F_M.MRAM\[29\]\[1\] _1539_ _1809_ mod.Data_Mem.F_M.MRAM\[28\]\[1\]
+ _2191_ _2192_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_2
X_4503_ _1173_ _1174_ _1175_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_117_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8271_ _0367_ net1 mod.Data_Mem.F_M.MRAM\[768\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__5118__A1 _1783_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5483_ _2096_ _2129_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_144_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5669__A2 _2118_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7222_ _3570_ _0333_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4434_ _1016_ _1021_ _1107_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_160_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_132_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7153_ _3242_ _3529_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_154_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4365_ _0948_ _1025_ _1038_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_113_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7124__S _3506_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_717 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6104_ _2718_ _2719_ _2720_ _2721_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_140_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_59_739 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7084_ mod.Data_Mem.F_M.MRAM\[21\]\[5\] _3489_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4296_ _0965_ _0969_ _0970_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_98_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_836 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_363 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6035_ _2539_ _2650_ _2652_ _2435_ _2653_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_100_335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6094__A2 mod.Data_Mem.F_M.MRAM\[790\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_858 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_74_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_396 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2208 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2219 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_66_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7986_ mod.Instr_Mem.instruction\[11\] net2 net1 mod.P1.instr_reg\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XPHY_14 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_54_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1507 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_25 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1518 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_36 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_54_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1529 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_1200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XPHY_47 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_54_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6937_ _3248_ _3399_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XPHY_58 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_35_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6868_ _3356_ _0193_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__8102__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5357__A1 mod.Data_Mem.F_M.MRAM\[799\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5819_ _2440_ _2441_ _2442_ _2443_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_167_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7593__I _3786_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6799_ _3315_ _3316_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_22_396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_536 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8538_ _0042_ net1 mod.Data_Mem.F_M.out_data\[34\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_108_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5109__A1 mod.Data_Mem.F_M.MRAM\[783\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8469_ _0565_ net1 mod.Data_Mem.F_M.MRAM\[796\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_163_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8252__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_1048 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8076__D mod.P3.Res\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6085__A2 _2201_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4096__A1 _0754_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_761 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_1111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2720 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_904 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2731 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2742 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2753 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2764 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_32_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_31 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2775 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2786 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2797 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_159_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5348__A1 _1700_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7209__S _3562_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4020__A1 mod.Arithmetic.CN.I_in\[23\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_1126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_114_427 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4323__A2 mod.Arithmetic.CN.I_in\[51\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5751__I _2375_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_801 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4150_ _0651_ mod.Arithmetic.CN.I_in\[33\] _0826_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_68_525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6068__B _1495_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6076__A2 _2692_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6783__S _3300_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4081_ _0728_ _0729_ _0758_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_49_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_1192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_110_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7840_ _0080_ _3171_ _3921_ _3916_ _3922_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_58_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6515__C _3118_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8125__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_145_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_51_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7771_ _3309_ mod.Data_Mem.F_M.MRAM\[797\]\[3\] _3878_ _3882_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__5587__B2 _2178_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4983_ _1561_ _1651_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_51_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6722_ _3264_ _0139_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_108_1020 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3934_ _0612_ _0080_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_108_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6653_ mod.Data_Mem.F_M.MRAM\[25\]\[6\] _3217_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_149_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6531__B _2394_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4830__I _1495_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5604_ mod.Data_Mem.F_M.MRAM\[29\]\[5\] _2226_ _2227_ mod.Data_Mem.F_M.MRAM\[28\]\[5\]
+ _2239_ _2240_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XANTENNA__8275__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4011__A1 _0687_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_722 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_20_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6584_ _3178_ _3179_ _3181_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__4011__B2 mod.Arithmetic.I_out\[73\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8323_ _0419_ net1 mod.Data_Mem.F_M.MRAM\[776\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_118_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5535_ _2167_ _2175_ _2176_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_106_917 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8254_ _0350_ net1 mod.Data_Mem.F_M.MRAM\[31\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5466_ _2111_ _2112_ _2114_ _2115_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_7205_ _3539_ mod.Data_Mem.F_M.MRAM\[29\]\[7\] _3549_ _3560_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4417_ mod.Arithmetic.CN.I_in\[36\] _1090_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5511__A1 _2152_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_114_950 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8185_ _0295_ net1 mod.Data_Mem.F_M.MRAM\[3\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5397_ _2058_ _0007_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5362__I1 mod.Data_Mem.F_M.MRAM\[0\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_503 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7136_ _3512_ _3518_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_4348_ _1004_ _1016_ _1021_ _1022_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_141_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7067_ _3480_ _0268_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4279_ _0687_ _0804_ _0953_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_41_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4078__B2 _0754_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6018_ _2352_ _2636_ _2354_ _2637_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_67_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2005 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2016 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_904 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2027 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2038 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1304 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2049 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1326 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7969_ _0195_ net1 mod.Data_Mem.F_M.MRAM\[6\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1337 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1359 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4941__S _1609_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4250__A1 _0637_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7319__A2 _3626_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_981 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6160__C _2775_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5750__A1 _1595_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_108_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_112_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5502__A1 _2143_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5353__I1 mod.Data_Mem.F_M.MRAM\[784\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5571__I _1548_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_609 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_104_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6058__A2 mod.Data_Mem.F_M.MRAM\[5\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_878 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8148__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3240 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8534__D _0038_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4915__I _1564_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3251 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3262 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_19_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2550 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5569__A1 _2184_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2561 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2572 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_745 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2583 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4851__S _1519_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_1130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2594 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8298__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1860 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4241__A1 _0915_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1871 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_20_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1882 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1893 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7030__I1 mod.Data_Mem.F_M.MRAM\[18\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_158_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5320_ _1967_ _1976_ _1977_ _1983_ _1984_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_127_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5251_ mod.Data_Mem.F_M.MRAM\[791\]\[4\] mod.Data_Mem.F_M.MRAM\[788\]\[4\] mod.Data_Mem.F_M.MRAM\[789\]\[4\]
+ mod.Data_Mem.F_M.MRAM\[790\]\[4\] _1829_ _1915_ _1916_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_47_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_114_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4202_ _0872_ _0874_ _0876_ _0877_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_151_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5182_ _1845_ mod.Data_Mem.F_M.MRAM\[773\]\[3\] _1847_ _1848_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_123_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7246__A1 _3294_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6049__A2 mod.Data_Mem.F_M.MRAM\[19\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4133_ _0808_ _0809_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_29_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_1129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6454__C1 _3060_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4064_ _0737_ _0740_ _0741_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_83_325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_83_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4825__I mod.Data_Mem.F_M.src\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_83_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7823_ _3171_ _3908_ _3912_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_64_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_169_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7754_ _3866_ _3872_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_24_469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_1203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4966_ _1620_ _1632_ _1633_ mod.Data_Mem.F_M.MRAM\[15\]\[1\] _1634_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_6705_ _3253_ mod.Data_Mem.F_M.MRAM\[28\]\[5\] _3250_ _3254_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_7685_ _3836_ _0530_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6261__B _2873_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5980__A1 _2343_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4897_ _1565_ _1566_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__7021__I1 mod.Data_Mem.F_M.MRAM\[18\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6636_ _3208_ _0109_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_22_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_138_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6688__S _3237_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6567_ _3003_ _3158_ _3160_ _3168_ _0079_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_164_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_8306_ _0402_ net1 mod.Data_Mem.F_M.MRAM\[774\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_105_202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5518_ _2158_ _2093_ _2159_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_156_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_106_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6498_ _2353_ _2318_ _2536_ _2556_ _3102_ _3103_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_65_1007 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7485__A1 _3634_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_1187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8237_ _0333_ net1 mod.Data_Mem.F_M.MRAM\[2\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_133_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5335__I1 _1995_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5449_ _1951_ mod.Data_Mem.F_M.MRAM\[799\]\[0\] _2098_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__4299__A1 _0716_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5496__B1 _2140_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4299__B2 _0709_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_160_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8168_ mod.Data_Mem.F_M.out_data\[78\] net2 net1 mod.Arithmetic.I_out\[78\] vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XFILLER_102_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7119_ _3252_ _3508_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_75_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8099_ mod.Data_Mem.F_M.out_data\[9\] net2 net1 mod.Arithmetic.CN.I_in\[9\] vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_101_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5343__S0 _1910_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6460__A2 _2490_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_90_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8440__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1101 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1112 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_27_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1123 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_151_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_42_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6212__A2 _1789_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_169_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1156 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1167 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4223__A1 _0656_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1178 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4074__I1 mod.Arithmetic.I_out\[73\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_575 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8590__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4774__A2 _1438_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_168_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_6_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_156_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5723__A1 _1932_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_128_81 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6279__A2 _1907_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6397__I _2429_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5326__I1 mod.Data_Mem.F_M.MRAM\[0\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_152_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_907 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_739 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_929 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_105_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_81_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6451__A2 mod.Data_Mem.F_M.MRAM\[769\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_168_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4462__A1 _0635_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_572 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3070 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3081 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3092 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_391 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2380 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4820_ mod.Data_Mem.F_M.src\[8\] _1489_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_2391 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_21_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_57_1091 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5962__A1 _2264_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1690 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4751_ _1203_ mod.Arithmetic.CN.I_in\[46\] _1208_ _1340_ _1421_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XANTENNA__7003__I1 mod.Data_Mem.F_M.MRAM\[17\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7470_ _3640_ mod.Data_Mem.F_M.MRAM\[780\]\[2\] _3707_ _3710_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4682_ mod.Arithmetic.CN.I_in\[61\] _1135_ _1353_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_159_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8196__RN net2 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6421_ _3016_ _3029_ _0072_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_128_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_127_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6352_ _2884_ _2961_ _2962_ _2895_ _1725_ _2963_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_115_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5190__A2 _1855_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5303_ mod.Data_Mem.F_M.MRAM\[15\]\[5\] _1599_ _1967_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__8313__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5317__I1 mod.Data_Mem.F_M.MRAM\[16\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6283_ mod.Data_Mem.F_M.MRAM\[789\]\[4\] mod.Data_Mem.F_M.MRAM\[791\]\[4\] mod.Data_Mem.F_M.MRAM\[790\]\[4\]
+ mod.Data_Mem.F_M.MRAM\[788\]\[4\] _2448_ _2383_ _2896_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_8022_ _0231_ net1 mod.Data_Mem.F_M.MRAM\[15\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_142_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5144__C _1557_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5234_ _1898_ _1628_ _1899_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_130_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_69_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5165_ _1608_ _1830_ _1614_ _1831_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__7132__S _3513_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8463__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_99_1114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4116_ _0792_ _0793_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_56_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5096_ _1761_ _1762_ _1565_ _1763_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_56_358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8120__RN net2 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4047_ mod.Arithmetic.CN.I_in\[12\] _0724_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_72_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_169_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6770__I net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7806_ _3901_ _0586_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_13_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7242__I1 mod.Data_Mem.F_M.MRAM\[30\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_206 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_217 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__4205__A1 _0878_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_24_277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5998_ _2464_ _2615_ _2616_ _2539_ _2617_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_71_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7737_ _3862_ _0556_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5953__A1 _2266_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4949_ _1577_ _1592_ _1599_ _1617_ _1618_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_130_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_137_113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_32_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7668_ mod.Data_Mem.F_M.MRAM\[791\]\[2\] _3828_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_138_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6619_ mod.Data_Mem.F_M.MRAM\[24\]\[5\] _3200_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_7599_ _3612_ _3789_ _3791_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_4_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_152_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_165_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5181__A2 _1846_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_1184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_48_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6418__C1 _2361_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6808__I1 _3322_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7630__A1 _3322_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8111__RN net2 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6433__A2 _3032_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_678 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_1023 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6197__A1 _1910_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5244__I0 mod.Data_Mem.F_M.MRAM\[771\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7980__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_169_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8336__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_157_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5172__A2 _1837_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_136_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5960__S _2283_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8486__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_124_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6121__A1 _2373_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_726 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_748 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_759 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_79_984 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_645 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8102__RN net2 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6424__A2 _2278_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6791__S _3300_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_604 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6970_ mod.Data_Mem.F_M.dest\[4\] _3372_ _3420_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_111_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_53_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5921_ _2097_ mod.Data_Mem.F_M.MRAM\[786\]\[4\] _2542_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_53_339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1037 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_34_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_1164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5852_ _1814_ _2475_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_61_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_1066 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_726 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_167_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4803_ _1444_ _1452_ _1472_ _1473_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XANTENNA__6283__S1 _2383_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4738__A2 _1209_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8571_ _0075_ net1 mod.Data_Mem.F_M.out_data\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__6983__I0 _3399_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5783_ _2406_ _2407_ _2408_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_7522_ _3729_ mod.Data_Mem.F_M.MRAM\[782\]\[6\] _3739_ _3742_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4734_ mod.Arithmetic.CN.I_in\[63\] _1403_ _1404_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__4043__C _0630_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8169__RN net2 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7453_ mod.Data_Mem.F_M.MRAM\[778\]\[3\] _3700_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4665_ mod.Arithmetic.CN.I_in\[46\] _1335_ _1336_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_134_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_147_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6404_ _3009_ _2389_ _2384_ _2503_ _3012_ _3013_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
X_7384_ _3665_ _0400_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4596_ mod.P2.Rout_reg\[0\] _0672_ _1267_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_66_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6966__S _3414_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6335_ _1635_ _2005_ _2946_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_116_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_726 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6112__A1 _2540_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_1168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6266_ _2869_ _2878_ _2879_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__4994__B _1531_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_153_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_88_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8005_ _0214_ net1 mod.Data_Mem.F_M.MRAM\[13\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5217_ _1530_ _1882_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_69_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6197_ _1910_ _1743_ _2812_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__4674__A1 _1234_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5148_ _1813_ _1814_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_57_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4285__I _0958_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5079_ _1518_ _1746_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__8209__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4426__A1 _0833_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_1220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7596__I _3786_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6179__A1 _1585_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8359__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6974__I0 _3386_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_157_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_153_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5154__A2 _1819_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8079__D mod.P3.Res\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_134_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__7151__I0 _3527_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6103__A1 _1764_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_856 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_121_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_48_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4665__A1 mod.Arithmetic.CN.I_in\[46\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_1071 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_36_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_47_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6406__A2 _2387_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_1006 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5614__B1 _1749_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_141_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_169_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8542__D _0046_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_575 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6343__C _1898_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_149_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5917__A1 _2506_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_31_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_141_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_606 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_89_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_1037 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4450_ _1009_ _1013_ _1123_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__7876__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4381_ _0957_ _0960_ _0961_ _1054_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_112_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6120_ _1505_ _1511_ _2736_ _1575_ _2733_ _2737_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_125_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_501 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6051_ _2352_ _2668_ _2354_ _2669_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5002_ _1669_ _1670_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_100_539 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_965 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4408__A1 _0716_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5605__B1 mod.Data_Mem.F_M.MRAM\[798\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_497 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_1139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_53_125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6953_ _3410_ _0224_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_93_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4959__A2 _1627_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5081__A1 _1745_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8501__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4833__I mod.Data_Mem.F_M.src\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5904_ _2211_ _2525_ _2526_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_53_169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6884_ _3364_ _0201_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_50_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5835_ mod.Data_Mem.F_M.MRAM\[14\]\[1\] mod.Data_Mem.F_M.MRAM\[15\]\[1\] _2452_ _2459_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__5908__A1 _2127_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6956__I0 _3395_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5759__I1 mod.Data_Mem.F_M.MRAM\[783\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5908__B2 _2527_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8554_ _0058_ net1 mod.Data_Mem.F_M.out_data\[18\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_50_898 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5384__A2 _2045_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5766_ _2388_ _2389_ _2390_ _2290_ _2376_ _2391_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
X_7505_ _3731_ mod.Data_Mem.F_M.MRAM\[781\]\[7\] _3726_ _3732_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4717_ _1279_ _1282_ _1387_ _1388_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
X_8485_ _0581_ net1 mod.Data_Mem.F_M.MRAM\[798\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__5664__I _1686_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_163_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5697_ _2256_ mod.Data_Mem.F_M.MRAM\[29\]\[5\] _2325_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_135_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7436_ _3691_ _0426_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_30_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_68_1208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4648_ _1306_ _1318_ _1319_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_151_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_146_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6696__S _3237_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7367_ mod.Data_Mem.F_M.MRAM\[773\]\[0\] _3657_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_122_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4579_ _1061_ _1251_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_89_501 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_157_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6318_ _2886_ _2926_ _2929_ _2930_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_89_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7298_ _3615_ mod.Data_Mem.F_M.MRAM\[768\]\[4\] _3606_ _3616_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_104_867 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtiny_user_project_17 io_oeb[6] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_104_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xtiny_user_project_28 io_oeb[17] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
X_6249_ _2850_ _2857_ _2862_ _2863_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_103_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xtiny_user_project_39 io_oeb[28] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XANTENNA__8031__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_18_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4944__S _1612_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2902 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7320__S _3623_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2913 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_946 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2924 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2935 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8181__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2946 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2957 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2968 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2979 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_13_501 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_164_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_111_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_40_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6947__I0 _3405_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_13_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6572__A1 _0612_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7899__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_1207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5574__I _1601_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6324__A1 _2134_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4886__A1 _1554_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_107_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7124__I0 _3462_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_81 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_92 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8537__D _0041_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_1049 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8524__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_751 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_497 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7052__A2 _3466_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5749__I _2373_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_607 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3950_ mod.P2.Rout_reg\[0\] mod.P2.Rout_reg\[1\] _0627_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_16_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_1213 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_1009 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5620_ _1940_ _2253_ _2254_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__6563__A1 mod.Data_Mem.F_M.MRAM\[780\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6563__B2 _3164_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_904 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5551_ _2186_ _2190_ _2191_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_145_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_117_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_571 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_4502_ _0613_ mod.Arithmetic.CN.I_in\[21\] mod.Arithmetic.CN.I_in\[20\] _1174_ vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__and3_1
X_8270_ _0366_ net1 mod.Data_Mem.F_M.MRAM\[768\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__6315__A1 _2872_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5482_ _2110_ _2127_ _2128_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_7221_ _3569_ mod.Data_Mem.F_M.MRAM\[2\]\[5\] _3567_ _3570_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4433_ _1004_ _1016_ _1105_ _1106_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_99_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4877__A1 _1536_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__8054__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7152_ _3528_ _0305_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4364_ _0976_ _1024_ _1037_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_99_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6103_ _1764_ _1589_ _2720_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_115_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_675 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_7083_ _3488_ _0276_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4295_ _0966_ _0968_ _0969_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_98_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6034_ _2549_ _2049_ _2651_ _2652_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_397 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_67_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_100_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2209 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7985_ mod.Instr_Mem.instruction\[10\] net2 net1 mod.P1.instr_reg\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XANTENNA__6264__B _2715_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_15 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__5054__A1 _1674_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_26 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1508 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1519 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6936_ _3398_ _0219_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XPHY_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_42_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_48 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_74_1212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_59 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__4801__A1 _1459_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_168_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6929__I0 _3393_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6867_ mod.Data_Mem.F_M.MRAM\[6\]\[1\] _3356_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_23_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_50_640 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5818_ _2283_ mod.Data_Mem.F_M.MRAM\[773\]\[1\] _2442_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_10_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6554__A1 _2548_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6798_ net8 _3315_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_50_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8537_ _0041_ net1 mod.Data_Mem.F_M.out_data\[33\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5749_ _2373_ _2374_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6306__A1 _2876_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5109__A2 _1775_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8468_ _0564_ net1 mod.Data_Mem.F_M.MRAM\[796\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_108_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7419_ mod.Data_Mem.F_M.MRAM\[776\]\[2\] _3683_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_135_277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8399_ _0495_ net1 mod.Data_Mem.F_M.MRAM\[786\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_123_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_150_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_951 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_1216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8547__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_77_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5293__A1 _1954_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_1082 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_92_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7050__S _3469_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2710 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2721 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2732 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2743 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2754 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2765 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2776 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_426 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2787 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2798 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_13_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6545__A1 _2611_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5348__A2 _2010_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6545__B2 _2211_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4556__B1 _1114_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_51_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__8077__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_154_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_1086 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7345__I0 _3645_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7225__S _3567_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5808__B1 _2427_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7914__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4080_ _0753_ _0755_ _0756_ _0757_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_62_1160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4087__A2 _0751_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5284__A1 _1551_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7770_ _3881_ _0570_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_17_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4982_ _1565_ _1649_ _1650_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_63_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6721_ mod.Data_Mem.F_M.MRAM\[10\]\[3\] _3264_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_3933_ mod.I_addr\[0\] _0612_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_60_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6652_ _3216_ _0117_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_108_1065 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__7584__I0 _3754_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6536__A1 _2474_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5603_ _2228_ _2238_ _2239_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_6583_ _3180_ _0084_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4011__A2 mod.Arithmetic.I_out\[74\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8322_ _0418_ net1 mod.Data_Mem.F_M.MRAM\[776\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_117_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5534_ _2158_ _2168_ _2174_ _2175_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_117_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8253_ _0349_ net1 mod.Data_Mem.F_M.MRAM\[31\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5465_ _2113_ _2066_ _2114_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_105_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4986__C _1653_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_160_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_133_748 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7204_ _3559_ _0326_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4416_ _0982_ _1088_ _1089_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_8184_ _0294_ net1 mod.Data_Mem.F_M.MRAM\[3\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__5511__A2 mod.Data_Mem.F_M.MRAM\[31\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5396_ _2038_ _2057_ _2058_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_87_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7135_ _3517_ _0299_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6974__S _3423_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4347_ _1018_ _1019_ _1020_ _1021_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_98_150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_526 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7066_ mod.Data_Mem.F_M.MRAM\[20\]\[4\] _3480_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_86_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_645 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_1058 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4278_ _0881_ _0884_ _0952_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__4078__A2 _0751_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5275__A1 _1931_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6472__B1 _2524_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6017_ _2061_ mod.Data_Mem.F_M.MRAM\[18\]\[6\] _2635_ _2636_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_86_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2006 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_540 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2017 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2028 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2039 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1305 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1316 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7968_ _0194_ net1 mod.Data_Mem.F_M.MRAM\[6\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_42_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1327 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_426 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1338 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1349 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6919_ _3385_ _0215_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_70_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7899_ _0125_ net1 mod.Data_Mem.F_M.MRAM\[27\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__4250__A2 _0922_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_168_13 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_50_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_51_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_167_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_161_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_156_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_10_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_163_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5852__I _1814_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7937__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_7_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5502__A2 _2145_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_151_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_1002 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5073__B _1562_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_1013 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_1182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_104_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_65 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5266__A1 mod.Data_Mem.F_M.MRAM\[799\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6463__B1 _3009_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6683__I _3236_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6463__C2 _3023_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3230 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3241 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3252 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3263 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_787 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2540 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2551 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_73_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2562 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2573 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2584 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2595 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1850 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1861 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4241__A2 mod.Arithmetic.ACTI.x\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1872 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_971 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_159_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1883 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1894 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_155_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5250_ _1914_ _1915_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_64_1200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4201_ _0803_ _0875_ _0876_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_5181_ _1647_ _1846_ _1847_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_25_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7246__A2 _3464_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4132_ _0807_ mod.Arithmetic.CN.I_in\[25\] _0808_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_110_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_96_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6454__B1 _3059_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6454__C2 _2477_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4063_ mod.Arithmetic.I_out\[78\] _0739_ _0703_ mod.Arithmetic.CN.I_in\[22\] _0740_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_2
XFILLER_68_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_497 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_1004 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7822_ mod.I_addr\[0\] _3169_ _3911_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_52_713 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8242__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5002__I _1669_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7753_ _3871_ _0563_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4965_ _1616_ _1633_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5937__I _2402_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4863__S0 _1527_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4841__I _1509_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6704_ _3252_ _3253_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_33_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6509__A1 _1491_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7684_ mod.Data_Mem.F_M.MRAM\[792\]\[2\] _3836_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4896_ _1564_ _1565_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_149_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_32_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_20_643 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6635_ mod.Data_Mem.F_M.MRAM\[26\]\[5\] _3208_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__8392__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3991__A1 _0660_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6566_ _1966_ _3162_ _3167_ _3168_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_106_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8305_ _0401_ net1 mod.Data_Mem.F_M.MRAM\[774\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_145_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5517_ _2157_ _2158_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_6497_ _3047_ _3101_ _3102_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_8236_ _0332_ net1 mod.Data_Mem.F_M.MRAM\[2\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_161_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_105_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7485__A2 _3371_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5448_ _2096_ _2097_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__5335__I2 _1996_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_1199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5496__A1 _2119_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4299__A2 _0816_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_154_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5496__B2 _2133_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8167_ mod.Data_Mem.F_M.out_data\[77\] net2 net1 mod.Arithmetic.I_out\[77\] vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_5379_ mod.Data_Mem.F_M.MRAM\[771\]\[7\] mod.Data_Mem.F_M.MRAM\[770\]\[7\] _1903_
+ _2041_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_102_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7118_ _3507_ _0292_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_87_643 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_943 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8098_ mod.Data_Mem.F_M.out_data\[8\] net2 net1 mod.Arithmetic.CN.I_in\[8\] vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_87_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_7049_ _3471_ _0259_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_86_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5343__S1 _1590_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_540 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_167_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_27_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1113 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1124 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1146 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1157 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1168 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1179 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_63_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_70_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3982__A1 _0635_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5723__A2 mod.Data_Mem.F_M.MRAM\[796\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_575 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_124_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_1157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_124_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5487__A1 _2072_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8115__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_643 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_751 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_93_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8545__D _0049_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6119__S _1782_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7302__I _3318_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8265__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5958__S _2161_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4462__A2 _1017_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3060 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_80_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3071 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3082 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3093 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2370 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2381 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2392 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5757__I _2381_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_1081 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1680 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4750_ _1374_ _1378_ _1419_ _1420_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__7539__I0 _3725_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1691 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_119_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4681_ _1225_ _0995_ _1231_ _1351_ _1352_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_144_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6420_ _2184_ _3025_ _3028_ _3029_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__5714__A2 _2150_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_1019 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6351_ _1994_ _1995_ _2044_ _2962_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_128_895 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5302_ _1965_ _1966_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_143_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_115_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6282_ _2881_ _2895_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_103_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8021_ _0230_ net1 mod.Data_Mem.F_M.MRAM\[15\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_88_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5233_ _1799_ _1898_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_130_526 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4150__A1 _0651_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5164_ mod.Data_Mem.F_M.MRAM\[787\]\[3\] mod.Data_Mem.F_M.MRAM\[786\]\[3\] _1829_
+ _1830_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_97_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6537__B _2698_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_773 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_57_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4115_ mod.Arithmetic.ACTI.x\[7\] _0676_ _0789_ mod.Arithmetic.ACTI.x\[6\] _0792_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_97_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5095_ mod.Data_Mem.F_M.MRAM\[773\]\[2\] mod.Data_Mem.F_M.MRAM\[772\]\[2\] _1746_
+ _1762_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_37_540 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4046_ _0707_ _0708_ _0717_ _0720_ _0721_ _0722_ _0723_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XANTENNA__5868__S _2152_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5650__A1 _2281_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7778__I0 _3782_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7805_ mod.Data_Mem.F_M.MRAM\[7\]\[2\] _3901_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XPHY_207 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_5997_ mod.Data_Mem.F_M.MRAM\[784\]\[6\] mod.Data_Mem.F_M.MRAM\[785\]\[6\] _2331_
+ _2616_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_52_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_229 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_80_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_1001 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7736_ mod.Data_Mem.F_M.MRAM\[795\]\[4\] _3862_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_24_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_429 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_1181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4948_ _1563_ _1605_ _1611_ _1615_ _1616_ _1617_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XANTENNA__5953__A2 mod.Data_Mem.F_M.MRAM\[14\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_1045 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_162_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_71_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7667_ _3827_ _0521_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_123_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4879_ _1494_ _1548_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_166_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6618_ _3199_ _0100_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_123_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_119_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5705__A2 _2142_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7598_ _1682_ _3789_ _3790_ _0489_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__8138__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6549_ _1966_ _3139_ _3141_ _3148_ _3151_ _0078_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai32_1
XFILLER_134_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_106_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5469__A1 _2116_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8219_ _0320_ net1 mod.Data_Mem.F_M.MRAM\[29\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__7831__B _3916_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_160_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6130__A2 _2200_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8288__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_1152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_1163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_751 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_1196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6418__B1 _2365_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6418__C2 _2672_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_784 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_540 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7630__A2 _3798_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5641__A1 _2063_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4444__A2 _1113_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_584 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7769__I0 _3306_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6197__A2 _1743_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_604 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_168_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_23_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_7_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4380__A1 _0617_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_1036 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_152_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_716 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7233__S _3574_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_738 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4132__A1 _0807_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_749 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5261__B _1925_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7032__I _3255_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_465 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5632__A1 _2264_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_1110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5920_ mod.Data_Mem.F_M.MRAM\[784\]\[4\] mod.Data_Mem.F_M.MRAM\[785\]\[4\] _2540_
+ _2541_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_46_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_146_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_1049 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_1045 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5851_ _1535_ _2474_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_62_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_1078 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4802_ _1454_ _1457_ _1471_ _1472_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XANTENNA__4199__A1 mod.Arithmetic.CN.I_in\[24\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8570_ _0074_ net1 mod.Data_Mem.F_M.out_data\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_21_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5782_ mod.Data_Mem.F_M.MRAM\[786\]\[0\] mod.Data_Mem.F_M.MRAM\[787\]\[0\] _1769_
+ _2407_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__6983__I1 mod.Data_Mem.F_M.MRAM\[16\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7521_ _3741_ _0461_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4733_ mod.Arithmetic.CN.I_in\[61\] _1366_ _1403_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_159_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_148_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7452_ _3699_ _0434_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4664_ _1202_ mod.Arithmetic.CN.I_in\[45\] _1335_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_107_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5699__A1 _2326_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6403_ _2422_ _3010_ _3011_ _3012_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_7383_ mod.Data_Mem.F_M.MRAM\[774\]\[0\] _3665_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4595_ _0799_ _0857_ _1266_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_128_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6111__I _1691_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6334_ _2870_ _2004_ _2945_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__8430__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6265_ _2871_ _2874_ _2875_ _2877_ _2878_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_142_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6112__A2 mod.Data_Mem.F_M.MRAM\[2\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8004_ _0213_ net1 mod.Data_Mem.F_M.MRAM\[13\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__4123__A1 _0661_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5216_ _1607_ _1881_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_69_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6196_ _1751_ _1747_ _2811_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_97_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_462 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4674__A2 _1344_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8580__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5147_ _1517_ _1813_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_56_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_84_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_977 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5078_ _1572_ _1745_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__4426__A2 _1097_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6781__I net4 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4029_ _0675_ _0705_ _0706_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_71_126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_13_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5397__I _2058_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6974__I1 mod.Data_Mem.F_M.MRAM\[16\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7719_ _3853_ _0547_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_138_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_165_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_158_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_109_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_107_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_106_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_162_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_106_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_45_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_69_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6103__A2 _1589_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7151__I1 mod.Data_Mem.F_M.MRAM\[12\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_161_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_121_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5081__B _1562_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4665__A2 _1335_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8095__D mod.Data_Mem.F_M.out_data\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_782 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_646 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5614__A1 mod.Data_Mem.F_M.MRAM\[797\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8096__RN net2 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6691__I _3242_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5614__B2 mod.Data_Mem.F_M.MRAM\[796\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_936 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_169_1157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_91_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8303__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5917__A2 mod.Data_Mem.F_M.MRAM\[788\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8453__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_157_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7027__I _3447_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5971__S _2540_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_1169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_651 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4380_ _0617_ _0680_ _0682_ _1053_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__5550__B1 _1632_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_153_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_124_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_846 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_513 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5153__I0 mod.Data_Mem.F_M.MRAM\[17\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_535 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6050_ _2129_ mod.Data_Mem.F_M.MRAM\[18\]\[7\] _2667_ _2668_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_546 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6087__B _2703_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_8509__189 net189 vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_112_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_568 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5001_ mod.Data_Mem.F_M.src\[8\] _1669_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_61_1033 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5853__A1 _2161_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_977 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4408__A2 _0816_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6952_ _3386_ mod.Data_Mem.F_M.MRAM\[15\]\[0\] _3409_ _3410_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_81_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5211__S _1875_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5081__A2 _1747_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5903_ _2517_ _2521_ _2523_ _2355_ _2524_ _2357_ _2525_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_1
X_6883_ mod.Data_Mem.F_M.MRAM\[4\]\[1\] _3364_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_50_800 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4335__B mod.Arithmetic.ACTI.x\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6106__I _1737_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5834_ mod.Data_Mem.F_M.MRAM\[30\]\[1\] _1632_ _2398_ _2458_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_22_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6956__I1 mod.Data_Mem.F_M.MRAM\[15\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6030__A1 _2428_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_1151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_1162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8553_ _0057_ net1 mod.Data_Mem.F_M.out_data\[17\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5765_ mod.Data_Mem.F_M.MRAM\[772\]\[0\] mod.Data_Mem.F_M.MRAM\[773\]\[0\] _1951_
+ _2390_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_72_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_1184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7504_ _3321_ _3731_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4592__A1 _0786_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4716_ _1324_ _1327_ _1386_ _1387_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
X_8484_ _0580_ net1 mod.Data_Mem.F_M.MRAM\[798\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5696_ _2324_ _0052_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_7435_ mod.Data_Mem.F_M.MRAM\[777\]\[2\] _3691_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_147_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4647_ _1174_ _1309_ _1317_ _1318_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
X_7366_ _3656_ _0391_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_144_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4578_ mod.Arithmetic.CN.I_in\[61\] _1250_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_116_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6776__I _3297_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6317_ _2718_ _2927_ _2928_ _2929_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_7297_ _3311_ _3615_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_1_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_143_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7970__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_879 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7833__A2 _3917_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6248_ _2108_ _2224_ _2861_ _2862_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
Xtiny_user_project_18 io_oeb[7] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_77_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xtiny_user_project_29 io_oeb[18] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XANTENNA__5844__A1 _2464_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_162_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_103_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6179_ _1585_ _2793_ _2794_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_131_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7601__S _3787_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8326__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8078__RN net2 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7597__A1 _3610_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2903 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_17_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_796 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2914 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2925 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2936 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_84_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6444__C _2073_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2947 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2958 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2969 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_513 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_1084 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8476__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6947__I1 mod.Data_Mem.F_M.MRAM\[14\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6021__A1 _2345_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7048__S _3469_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6572__A2 _3169_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_139_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_153_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_426 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6324__A2 mod.Data_Mem.F_M.MRAM\[15\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4335__A1 mod.Arithmetic.CN.I_in\[64\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5383__I0 _2040_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_651 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_1180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4886__A2 _1537_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6686__I net4 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5590__I _1600_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7124__I1 mod.Data_Mem.F_M.MRAM\[3\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6088__A1 _2012_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7824__A2 _3911_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7511__S _3734_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_966 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_977 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_796 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8553__D _0057_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_690 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_1157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_1037 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_31_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6563__A2 _1674_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5550_ _2188_ mod.Data_Mem.F_M.MRAM\[30\]\[1\] _1632_ _2189_ _2190_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
X_4501_ _0678_ mod.Arithmetic.CN.I_in\[20\] _0843_ _1173_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_129_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5481_ mod.Data_Mem.F_M.MRAM\[30\]\[3\] mod.Data_Mem.F_M.MRAM\[31\]\[3\] _1845_ _2127_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__6315__A2 _1958_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7220_ _3252_ _3569_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4326__A1 _0993_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5374__I0 _2032_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4432_ _1018_ _1020_ _1104_ _1105_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_126_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7993__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_67_1220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7151_ _3527_ mod.Data_Mem.F_M.MRAM\[12\]\[1\] _3525_ _3528_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4363_ _0861_ _0938_ _1027_ _1036_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_98_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_154_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6102_ _2186_ _1582_ _2719_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_99_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7082_ mod.Data_Mem.F_M.MRAM\[21\]\[4\] _3488_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4294_ _0868_ _0966_ _0967_ _0968_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_86_505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8349__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_101_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6033_ _2097_ mod.Data_Mem.F_M.MRAM\[786\]\[7\] _2651_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_398 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_67_752 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_711 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6037__S _2326_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7220__I _3252_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8499__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7984_ mod.Instr_Mem.instruction\[9\] net2 net1 mod.P1.instr_reg\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XANTENNA__6251__A1 _2079_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_16 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1509 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_27 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_6935_ _3397_ mod.Data_Mem.F_M.MRAM\[14\]\[3\] _3391_ _3398_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XPHY_38 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_81_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_49 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__4801__A2 _1463_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6929__I1 mod.Data_Mem.F_M.MRAM\[14\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6866_ _3355_ _0192_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6003__A1 _2619_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5817_ _2281_ mod.Data_Mem.F_M.MRAM\[772\]\[1\] _2441_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6797_ _3314_ _0164_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6554__A2 _2673_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4565__A1 _1124_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8536_ _0040_ net1 mod.Data_Mem.F_M.out_data\[32\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5748_ _1542_ _1533_ _2373_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_109_916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_927 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_426 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6306__A2 _1973_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8467_ _0563_ net1 mod.Data_Mem.F_M.MRAM\[796\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5679_ _2089_ _2131_ _2307_ _2308_ _2309_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_68_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4317__A1 _0921_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_151_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7418_ _3682_ _0417_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5365__I0 mod.Data_Mem.F_M.MRAM\[5\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8398_ _0494_ net1 mod.Data_Mem.F_M.MRAM\[786\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_117_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_610 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7349_ _3620_ mod.Data_Mem.F_M.MRAM\[771\]\[7\] _3643_ _3648_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_89_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_974 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5817__A1 _2281_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_1050 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_77_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7331__S _3636_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5293__A2 _1955_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_1113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_936 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2700 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2711 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_17_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2722 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2733 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2744 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2755 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7866__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2766 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2777 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2788 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2799 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4703__B _0634_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6545__A2 _2627_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4556__A1 _0645_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_166_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7345__I1 mod.Data_Mem.F_M.MRAM\[771\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4308__A1 _0980_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_147_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_971 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_154_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_135_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7305__I _3321_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_110_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5808__A1 _2423_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_836 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5808__B2 _2403_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_730 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5284__A2 _1939_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6481__A1 _2264_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6365__B _2715_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_76_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7040__I _3465_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6084__C _1965_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6233__A1 _1802_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4981_ mod.Data_Mem.F_M.MRAM\[1\]\[1\] mod.Data_Mem.F_M.MRAM\[0\]\[1\] _1509_ _1649_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_51_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6720_ _3263_ _0138_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA_output6_I net6 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_147_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7033__I0 _3460_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6651_ mod.Data_Mem.F_M.MRAM\[25\]\[5\] _3216_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_5602_ _1953_ mod.Data_Mem.F_M.MRAM\[31\]\[5\] mod.Data_Mem.F_M.MRAM\[30\]\[5\] _2229_
+ _2238_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XANTENNA__8021__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4547__A1 _1205_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6582_ _3178_ _3179_ _3180_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_164_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_158_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8321_ _0417_ net1 mod.Data_Mem.F_M.MRAM\[776\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5533_ mod.Data_Mem.F_M.MRAM\[797\]\[0\] _1729_ _2173_ _2174_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_8_380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_117_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8252_ _0348_ net1 mod.Data_Mem.F_M.MRAM\[31\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_133_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5464_ _1803_ _2113_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_7203_ _3537_ mod.Data_Mem.F_M.MRAM\[29\]\[6\] _3553_ _3559_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__8171__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4415_ _0986_ _1088_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_8183_ _0293_ net1 mod.Data_Mem.F_M.MRAM\[3\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_126_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5395_ _2039_ _2046_ _2056_ _1927_ _1629_ _2057_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_99_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7134_ _3454_ mod.Data_Mem.F_M.MRAM\[19\]\[3\] _3513_ _3517_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_154_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4346_ _0813_ _0923_ _0840_ _1020_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_98_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_674 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6847__I0 _3259_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7065_ _3479_ _0267_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_59_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4277_ _0947_ _0949_ _0935_ _0950_ _0889_ _0951_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai32_1
XFILLER_98_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7151__S _3525_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6472__A1 _3021_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6016_ _1685_ mod.Data_Mem.F_M.MRAM\[19\]\[6\] _2635_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__5275__A2 _1936_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6472__B2 _3009_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7889__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_55_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2007 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2018 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6224__A1 _1931_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2029 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1306 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_7967_ _0193_ net1 mod.Data_Mem.F_M.MRAM\[6\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_55_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1317 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1328 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1339 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4786__A1 mod.Arithmetic.CN.I_in\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_78_1190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6918_ _3259_ mod.Data_Mem.F_M.MRAM\[13\]\[7\] _3381_ _3385_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_70_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_168_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7898_ _0124_ net1 mod.Data_Mem.F_M.MRAM\[27\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_23_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7024__I0 _3454_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_1054 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6849_ mod.Data_Mem.F_M.MRAM\[779\]\[0\] _3347_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_23_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6527__A2 _3130_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4538__A1 mod.Arithmetic.CN.I_in\[43\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8519_ net183 net1 mod.Data_Mem.F_M.out_data\[63\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__8514__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_746 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_148_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7326__S _3625_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_501 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_108_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4710__A1 _1372_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_117_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_78_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_1194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5266__A2 _1599_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6463__A1 _3005_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6463__B2 _2487_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_18_402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_711 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3220 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3231 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3242 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3253 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6215__A1 _1800_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7263__I0 mod.Data_Mem.F_M.MRAM\[31\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2530 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2541 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2552 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2563 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2574 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8044__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4777__A1 _1297_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1840 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2585 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2596 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1851 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7015__I0 _3445_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1862 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_158_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1873 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1884 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_1127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_92_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6518__A2 _3121_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1895 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_105_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_146_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8194__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4659__I mod.Arithmetic.CN.I_in\[37\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7035__I _3258_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_1212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4200_ _0844_ mod.Arithmetic.CN.I_in\[18\] _0875_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_69_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5180_ mod.Data_Mem.F_M.MRAM\[772\]\[3\] _1846_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_111_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_111_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4131_ _0806_ _0807_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_96_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7246__A3 _3296_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_111_966 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6454__A1 _2503_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6454__B2 _2568_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_465 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4062_ _0738_ _0739_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_83_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6206__A1 _1730_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7821_ _3910_ _0592_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_92_872 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_393 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7752_ _3309_ mod.Data_Mem.F_M.MRAM\[796\]\[3\] _3867_ _3871_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4964_ mod.Data_Mem.F_M.MRAM\[31\]\[1\] _1632_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4863__S1 _1531_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6703_ net8 _3252_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_71_1216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8537__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7683_ _3835_ _0529_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4895_ _1525_ _1564_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_32_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6634_ _3207_ _0108_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__3991__A2 _0667_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_165_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5193__A1 _1642_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6565_ _3017_ _3163_ _3165_ _3166_ _3167_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_118_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8304_ _0400_ net1 mod.Data_Mem.F_M.MRAM\[774\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5516_ _1543_ _2157_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_106_716 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6496_ _2103_ _2559_ _3101_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_105_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_1167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_160_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_8235_ _0331_ net1 mod.Data_Mem.F_M.MRAM\[2\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_105_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6985__S _3428_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5447_ _1522_ _2096_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5335__I3 _1997_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5496__A2 _2137_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5740__I0 mod.Data_Mem.F_M.MRAM\[18\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5378_ mod.Data_Mem.F_M.MRAM\[769\]\[7\] mod.Data_Mem.F_M.MRAM\[768\]\[7\] _1814_
+ _2040_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_8166_ mod.Data_Mem.F_M.out_data\[76\] net2 net1 mod.Arithmetic.I_out\[76\] vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_99_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7117_ _3456_ mod.Data_Mem.F_M.MRAM\[3\]\[4\] _3506_ _3507_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4329_ _0913_ _0920_ _1003_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_87_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8097_ mod.Data_Mem.F_M.out_data\[7\] net2 net1 mod.Arithmetic.ACTI.x\[7\] vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_59_335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7493__I0 _3711_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_817 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7048_ _3454_ mod.Data_Mem.F_M.MRAM\[1\]\[3\] _3469_ _3471_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_87_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_101_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_722 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8067__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7829__B _3908_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_500 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_15_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1103 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1114 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1125 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1136 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1158 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1169 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_137_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7904__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3982__A2 mod.Arithmetic.CN.I_in\[56\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5184__A1 _1614_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_155_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7056__S _3465_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_1212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_152_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_21 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_100_1169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_151_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_105_771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_78_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6694__I net6 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_730 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_104_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6436__A1 _2071_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_891 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4998__A1 _1664_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3050 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4462__A3 _1134_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_3061 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3072 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3083 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_894 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3094 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_34_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8561__D _0065_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2360 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2371 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2382 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2393 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_159_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1681 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7539__I1 _1901_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1692 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_105_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_1014 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4680_ _1227_ _1230_ _1351_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_41_290 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_147_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6869__I mod.Data_Mem.F_M.MRAM\[6\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5773__I _1658_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6350_ _1997_ _1996_ _1713_ _2961_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__4922__A1 _1585_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5301_ _1964_ _1965_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_52_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__4389__I mod.Arithmetic.CN.I_in\[28\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6281_ _2886_ _2889_ _2893_ _2894_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_115_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8020_ _0229_ net1 mod.Data_Mem.F_M.MRAM\[15\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__6675__A1 mod.Data_Mem.F_M.dest\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5232_ _1888_ _1896_ _1633_ _1897_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_64_1020 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5163_ _1816_ _1829_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__4150__A2 mod.Arithmetic.CN.I_in\[33\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_430 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6427__A1 _2728_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_975 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4114_ _0783_ _0787_ _0790_ _0791_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_69_677 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_96_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_151_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5094_ mod.Data_Mem.F_M.MRAM\[775\]\[2\] mod.Data_Mem.F_M.MRAM\[774\]\[2\] _1746_
+ _1761_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_57_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4989__A1 _1655_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4045_ mod.Arithmetic.CN.I_in\[11\] _0722_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XANTENNA__5013__I _1676_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5650__A2 mod.Data_Mem.F_M.MRAM\[29\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_574 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6553__B _2381_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_894 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7778__I1 mod.Data_Mem.F_M.MRAM\[797\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4852__I mod.Data_Mem.F_M.src\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7804_ _3900_ _0585_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6045__S _2540_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7927__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_52_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_219 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_24_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5996_ _2313_ _2013_ _2614_ _2615_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__6272__C _1490_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_12_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7735_ _3861_ _0555_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_52_588 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4947_ _1506_ _1616_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_40_739 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_1193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_36_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7666_ mod.Data_Mem.F_M.MRAM\[791\]\[1\] _3827_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4878_ _1508_ _1532_ _1533_ _1546_ _1547_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_20_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6617_ mod.Data_Mem.F_M.MRAM\[24\]\[4\] _3199_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_137_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5683__I _2311_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7597_ _3610_ _3789_ _3790_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_118_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6548_ _1491_ _3150_ _3151_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_161_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6479_ _3083_ _1855_ _3084_ _3085_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_121_505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8218_ _0319_ net1 mod.Data_Mem.F_M.MRAM\[22\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_134_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4141__A2 _0816_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8149_ mod.Data_Mem.F_M.out_data\[59\] net2 net1 mod.Arithmetic.CN.I_in\[59\] vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_88_975 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6418__A1 _3026_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7466__I0 _3603_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6418__B2 _3006_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_796 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7218__I0 _3533_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_393 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_169_785 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_157_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_15_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5157__A1 _1653_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5807__B _2429_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6354__B1 mod.Data_Mem.F_M.MRAM\[14\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_1091 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4380__A2 _0680_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8232__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4002__I _0678_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_1048 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_48_1059 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_155_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_717 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5865__C1 _2487_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_739 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_430 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_97_249 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7313__I _3625_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5034__S _1701_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6409__A1 _2171_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8382__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7209__I0 _3523_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5632__A2 mod.Data_Mem.F_M.MRAM\[29\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1017 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_93_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_820 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_1144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5850_ _2467_ _2472_ _2473_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_94_1057 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2190 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4801_ _1459_ _1463_ _1470_ _1471_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XANTENNA__4199__A2 _0809_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5781_ _2109_ _2406_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_7520_ _3645_ mod.Data_Mem.F_M.MRAM\[782\]\[5\] _3739_ _3741_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4732_ _1400_ _1384_ _1401_ _1402_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_9_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_7451_ mod.Data_Mem.F_M.MRAM\[778\]\[2\] _3699_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4663_ mod.Arithmetic.CN.I_in\[38\] _1332_ _1333_ _1334_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_119_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5209__S _1873_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5699__A2 mod.Data_Mem.F_M.MRAM\[28\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6402_ _2256_ mod.Data_Mem.F_M.MRAM\[781\]\[0\] _3011_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_7382_ _3664_ _0399_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4594_ _1031_ _1262_ _1264_ _1265_ mod.P3.Res\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_6333_ _2866_ _2944_ _0069_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_143_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_66_1126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_115_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6499__I1 mod.Data_Mem.F_M.MRAM\[782\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_6264_ _2876_ _1878_ _2715_ _2877_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_131_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8003_ _0212_ net1 mod.Data_Mem.F_M.MRAM\[13\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5215_ mod.Data_Mem.F_M.MRAM\[3\]\[4\] mod.Data_Mem.F_M.MRAM\[2\]\[4\] _1879_ _1880_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_6195_ _2759_ _2806_ _2809_ _2810_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_85_901 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5146_ _1811_ _1812_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_97_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5879__S _2161_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5077_ _1742_ _1743_ _1744_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_38_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4028_ _0674_ mod.Arithmetic.I_out\[79\] _0705_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_56_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_820 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_680 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_80_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_1108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8105__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_536 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5979_ _2301_ mod.Data_Mem.F_M.MRAM\[773\]\[5\] _2599_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_7718_ mod.Data_Mem.F_M.MRAM\[794\]\[3\] _3853_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_139_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_166_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5627__B _2259_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7649_ _3818_ _0512_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_20_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_60_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__8255__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_800 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_1204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7334__S _3636_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_47_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_87_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_102_571 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_76_945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_1019 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7509__S _3734_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6413__S _2258_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_1090 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_169_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6327__B1 mod.Data_Mem.F_M.MRAM\[782\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_1096 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_1104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5925__I0 mod.Data_Mem.F_M.MRAM\[782\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_125_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5550__A1 _2188_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5550__B2 _2189_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7244__S _3579_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_152_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_503 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_525 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4667__I mod.Arithmetic.CN.I_in\[45\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4105__A2 _0774_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5153__I1 mod.Data_Mem.F_M.MRAM\[16\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_536 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6350__I0 _1997_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_1181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_761 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5000_ _1654_ _1667_ _1622_ _1668_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_569 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_1023 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_1045 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_113_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_93_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5605__A2 mod.Data_Mem.F_M.MRAM\[799\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_617 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_96_1119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_53_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6951_ _3408_ _3409_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__8128__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5902_ mod.Data_Mem.F_M.MRAM\[2\]\[3\] mod.Data_Mem.F_M.MRAM\[3\]\[3\] _2321_ _2524_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_81_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6882_ _3363_ _0200_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4335__C _0643_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_981 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5369__A1 mod.Data_Mem.F_M.MRAM\[31\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5833_ _2366_ _2457_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_61_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_536 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8278__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_569 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8552_ _0056_ net1 mod.Data_Mem.F_M.out_data\[16\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_72_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5764_ mod.Data_Mem.F_M.MRAM\[770\]\[0\] mod.Data_Mem.F_M.MRAM\[771\]\[0\] _1581_
+ _2389_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_50_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_148_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7503_ _3730_ _0454_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4715_ _1347_ _1385_ _1386_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_8483_ _0579_ net1 mod.Data_Mem.F_M.MRAM\[798\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_72_1196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5695_ _2082_ _2318_ _2323_ _2306_ _2324_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__6122__I _2706_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7434_ _3690_ _0425_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4646_ _1312_ _1316_ _1317_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_116_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5541__A1 _1782_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7365_ mod.Data_Mem.F_M.MRAM\[772\]\[7\] _3656_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4577_ _1240_ _1248_ _1249_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__7154__S _3525_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5541__B2 _2009_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6316_ _2891_ _1957_ _2928_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_131_611 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7296_ _1855_ _3609_ _3614_ _0363_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_103_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7294__A1 _1770_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6341__I0 mod.Data_Mem.F_M.MRAM\[789\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6247_ _2107_ _2860_ _2202_ _2210_ _2861_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_44_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xtiny_user_project_19 io_oeb[8] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_103_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5844__A2 _2466_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6178_ _2319_ mod.Data_Mem.F_M.MRAM\[783\]\[2\] mod.Data_Mem.F_M.MRAM\[782\]\[2\]
+ _2311_ _2793_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_97_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5910__B _2531_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5129_ _1781_ _1786_ _1789_ _1794_ _1527_ _1795_ _1796_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_57_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_606 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2904 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2915 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2926 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2937 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2948 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2959 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_129_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4280__A1 _0871_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6021__A2 mod.Data_Mem.F_M.MRAM\[4\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_878 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5080__I0 mod.Data_Mem.F_M.MRAM\[19\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6460__C _3047_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5357__B _2019_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5780__A1 _2403_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5907__I0 mod.Data_Mem.F_M.MRAM\[16\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_154_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_107_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5532__A1 _2169_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5383__I1 _2041_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_1192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_101_1094 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6188__B _2703_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_1007 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6088__A2 _1610_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_462 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_48_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8508__190 net190 vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_75_252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5599__A1 _1574_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_745 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8420__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_171 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_71_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4950__I _1499_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_1169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_1049 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_878 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_32_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4023__A1 _0696_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8570__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7038__I _3234_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5982__S _2522_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_157_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4500_ _1170_ _1171_ _1172_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_5480_ _1803_ _2126_ _0034_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4431_ _0824_ _1018_ _1020_ _1104_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__4326__A2 _0999_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7150_ _3239_ _3527_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4362_ _0945_ _1026_ _1035_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_99_823 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6101_ _2707_ _2718_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_7081_ _3487_ _0275_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_59_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4293_ _0878_ _0879_ _0870_ _0967_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_140_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_113_677 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_344 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_355 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6032_ mod.Data_Mem.F_M.MRAM\[784\]\[7\] mod.Data_Mem.F_M.MRAM\[785\]\[7\] _2331_
+ _2650_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_112_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_67_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_27_606 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7501__I _3318_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6545__C _3147_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_572 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7983_ mod.Instr_Mem.instruction\[8\] net2 net1 mod.P1.instr_reg\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_55_959 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_285 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_148_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_17 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_54_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6934_ _3245_ _3397_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XPHY_28 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_81_255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_39 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_63_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6865_ mod.Data_Mem.F_M.MRAM\[6\]\[0\] _3355_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_62_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_161_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6003__A2 mod.Data_Mem.F_M.MRAM\[782\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_161_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5816_ _2396_ _2440_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6796_ mod.Data_Mem.F_M.MRAM\[799\]\[4\] _3312_ _3313_ _3314_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_10_539 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8535_ _0039_ net1 mod.Data_Mem.F_M.out_data\[47\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5747_ _2353_ _2363_ _2371_ _1498_ _2372_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XANTENNA__5762__A1 _2385_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4565__A2 _1132_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7991__RN net2 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8466_ _0562_ net1 mod.Data_Mem.F_M.MRAM\[796\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5678_ _2295_ mod.Data_Mem.F_M.MRAM\[796\]\[3\] _2259_ _2308_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_136_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_159_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7417_ mod.Data_Mem.F_M.MRAM\[776\]\[1\] _3682_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5514__A1 _2138_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_1018 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5365__I1 mod.Data_Mem.F_M.MRAM\[4\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4629_ _1166_ _1298_ _1299_ _1300_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_8397_ _0493_ net1 mod.Data_Mem.F_M.MRAM\[786\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_116_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7348_ _3647_ _0382_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_1_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_131_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7279_ mod.Data_Mem.F_M.MRAM\[5\]\[7\] _3602_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_77_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5817__A2 mod.Data_Mem.F_M.MRAM\[772\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_539 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8443__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6455__C _3014_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2701 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2712 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2723 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2734 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_167_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2745 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_23 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2756 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2767 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_32_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2778 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2789 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8593__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4703__C mod.Arithmetic.ACTI.x\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4556__A2 mod.Arithmetic.CN.I_in\[53\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_1071 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_1033 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7982__RN net2 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5505__A1 _2135_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput3 net3 io_out[16] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XFILLER_108_994 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7522__S _3739_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4010__I _0682_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5808__A2 _2122_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_163_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8564__D _0068_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4945__I _1561_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5284__A3 _1947_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_1184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4492__A1 _1075_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_285 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_63_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_91_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6233__A2 _1832_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4980_ mod.Data_Mem.F_M.MRAM\[3\]\[1\] mod.Data_Mem.F_M.MRAM\[2\]\[1\] _1647_ _1648_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_52_929 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_981 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7033__I1 mod.Data_Mem.F_M.MRAM\[18\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_962 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6650_ _3215_ _0116_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_108_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7960__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6536__A3 _3138_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_995 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5601_ _2225_ _2232_ _2237_ _2178_ _0044_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_82_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6581_ _3175_ _3176_ _3179_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_31_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8320_ _0416_ net1 mod.Data_Mem.F_M.MRAM\[776\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_121_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_714 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5532_ _2169_ _2172_ _2173_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_118_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8316__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8251_ _0347_ net1 mod.Data_Mem.F_M.MRAM\[31\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5463_ mod.Data_Mem.F_M.MRAM\[30\]\[0\] mod.Data_Mem.F_M.MRAM\[31\]\[0\] _1873_ _2112_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_105_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7202_ _3558_ _0325_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6400__I _2499_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4414_ _0992_ _1085_ _1086_ _1023_ _0988_ _0989_ _1087_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai33_1
X_8182_ _0292_ net1 mod.Data_Mem.F_M.MRAM\[3\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5394_ mod.Data_Mem.F_M.MRAM\[799\]\[7\] _1913_ _2055_ _2056_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_7133_ _3516_ _0298_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_28_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4345_ _0617_ _1017_ _1019_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_114_975 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8466__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6847__I1 mod.Data_Mem.F_M.MRAM\[769\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7064_ mod.Data_Mem.F_M.MRAM\[20\]\[3\] _3479_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4276_ _0903_ _0934_ _0950_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_86_325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_859 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8150__RN net2 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6015_ _2548_ _2632_ _2633_ _2634_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_86_358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6472__A2 _2527_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2008 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2019 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6224__A2 _1817_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7966_ _0192_ net1 mod.Data_Mem.F_M.MRAM\[6\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1307 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1318 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_14_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_39_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1329 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6917_ _3384_ _0214_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_23_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5983__A1 _2398_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7897_ _0123_ net1 mod.Data_Mem.F_M.MRAM\[27\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__7024__I1 mod.Data_Mem.F_M.MRAM\[18\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6848_ _3346_ _0183_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_52_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_168_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_23_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_168_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4538__A2 _1096_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6779_ mod.Data_Mem.F_M.MRAM\[799\]\[0\] _3293_ _3300_ _3301_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__7607__S _3786_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8518_ net184 net1 mod.Data_Mem.F_M.out_data\[62\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_6_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8449_ _0545_ net1 mod.Data_Mem.F_M.MRAM\[794\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__3934__I _0612_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_164_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4031__S _0703_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_513 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_85_1162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4710__A2 _1380_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_986 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7342__S _3643_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_120_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_77_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6463__A2 _2298_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8141__RN net2 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3210 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3221 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_133_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3232 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_391 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3243 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3254 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6215__A2 _2818_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2520 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7263__I1 _3322_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2531 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2542 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7983__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2553 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2564 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2575 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5974__A1 _2410_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1830 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2586 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5596__I _1594_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1841 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2597 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1852 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_951 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1863 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7015__I1 mod.Data_Mem.F_M.MRAM\[18\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_13_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1874 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_984 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1885 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1896 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_1188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__8339__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_158_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4005__I mod.Arithmetic.CN.I_in\[18\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5037__S _1704_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8489__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_154_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6151__A1 _2180_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_290 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7252__S _3585_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4130_ mod.Arithmetic.CN.F_in\[0\] _0806_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_111_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_68_325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_859 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4061_ _0674_ _0677_ _0694_ _0700_ _0738_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XANTENNA__8132__RN net2 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6454__A2 _2478_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4465__A1 _0923_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_49_572 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_1093 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6206__A2 _1767_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7820_ _3907_ _3908_ _3909_ _3910_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_58_1006 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7254__I1 _3555_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_575 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4217__A1 _0891_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7751_ _3870_ _0562_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_52_759 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5965__A1 _1627_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4963_ _1628_ _1631_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6702_ _3251_ _0132_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_7682_ mod.Data_Mem.F_M.MRAM\[792\]\[1\] _3835_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4894_ _1562_ _1563_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_60_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6633_ mod.Data_Mem.F_M.MRAM\[26\]\[4\] _3207_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__8199__RN net2 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_164_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_678 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6564_ _2503_ _2655_ _2656_ _3050_ _3166_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_8303_ _0399_ net1 mod.Data_Mem.F_M.MRAM\[773\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5515_ _2119_ _2154_ _2156_ _2133_ _0039_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_121_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6495_ _2353_ _3095_ _3099_ _2108_ _3100_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_69_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8234_ _0330_ net1 mod.Data_Mem.F_M.MRAM\[2\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5446_ _2091_ _2094_ _2095_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__6142__A1 _2703_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_1179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8165_ mod.Data_Mem.F_M.out_data\[75\] net2 net1 mod.Arithmetic.I_out\[75\] vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XANTENNA__5740__I1 mod.Data_Mem.F_M.MRAM\[19\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5377_ mod.Data_Mem.F_M.MRAM\[783\]\[7\] _1673_ _2039_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_87_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7116_ _3500_ _3506_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_59_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5328__S0 _1881_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4328_ _1000_ _1001_ _1002_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_8096_ mod.Data_Mem.F_M.out_data\[6\] net2 net1 mod.Arithmetic.ACTI.x\[6\] vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_59_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8123__RN net2 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7047_ _3470_ _0258_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4259_ _0907_ _0927_ _0933_ _0934_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_74_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_68_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_167_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4208__A1 mod.Arithmetic.CN.I_in\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1104 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_15_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1126 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1137 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5956__A1 _2531_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7949_ _0175_ net1 mod.Data_Mem.F_M.MRAM\[789\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_70_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_169_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1148 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_63_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1159 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5708__A1 _2313_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7337__S _3636_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4392__B1 _1064_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7136__I _3512_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6133__A1 _2682_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_33 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_152_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_78_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_78_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8114__RN net2 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8011__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3040 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3051 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3062 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3073 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_3084 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3095 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2350 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2361 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8161__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2372 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2383 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2394 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5259__C _1642_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1660 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1671 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1682 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1693 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_146_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_159_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_105_1059 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7879__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_864 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4922__A2 _1589_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5300_ _1724_ _1964_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__6124__A1 _2738_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6280_ _2718_ _2890_ _2892_ _2893_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__6675__A2 mod.Data_Mem.F_M.dest\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5231_ _1889_ _1891_ _1893_ _1895_ _1751_ _1882_ _1896_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_103_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4686__A1 _0636_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_1054 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5162_ _1826_ _1827_ _1828_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_111_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_645 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8105__RN net2 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7624__A1 _1919_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4113_ _0786_ _0785_ _0789_ mod.Arithmetic.ACTI.x\[6\] _0790_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_57_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5093_ _1755_ _1758_ _1759_ _1760_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_97_987 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_1106 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_615 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4438__A1 _1109_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_1019 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_110_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4044_ _0680_ mod.Arithmetic.I_out\[75\] _0713_ _0721_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__4989__A2 _1656_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8504__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5230__S _1894_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7803_ mod.Data_Mem.F_M.MRAM\[7\]\[1\] _3900_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_52_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_5995_ _2214_ mod.Data_Mem.F_M.MRAM\[786\]\[6\] _2614_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_24_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7734_ mod.Data_Mem.F_M.MRAM\[795\]\[3\] _3861_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_24_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4946_ _1603_ _1613_ _1614_ _1615_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_7665_ _3826_ _0520_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4877_ _1536_ _1545_ _1546_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__7157__S _3525_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_165_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6616_ _3198_ _0099_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_20_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7596_ _3786_ _3789_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6996__S _3435_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6547_ _3111_ _3149_ _3150_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_152_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_106_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_536 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7163__I0 _3508_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6478_ _2315_ mod.Data_Mem.F_M.MRAM\[769\]\[3\] _3084_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_133_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_106_569 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8217_ _0318_ net1 mod.Data_Mem.F_M.MRAM\[22\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_134_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5429_ _1725_ _2084_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__8034__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_943 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8148_ mod.Data_Mem.F_M.out_data\[58\] net2 net1 mod.Arithmetic.CN.I_in\[58\] vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_0_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_82_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_753 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_58_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_59_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6418__A2 _2272_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8079_ mod.P3.Res\[7\] net2 net1 net10 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XANTENNA__7620__S _3801_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4429__A1 _1095_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8184__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7218__I1 mod.Data_Mem.F_M.MRAM\[2\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5140__S _1510_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_575 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_895 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5929__A1 _2549_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_167_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_1015 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_71_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4601__A1 _1149_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_169_797 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_11_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5157__A2 _1815_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6354__A1 _2134_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6354__B2 _2216_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7154__I0 _3529_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4380__A3 _0682_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_98_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4668__A1 _1203_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_718 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5315__S _1968_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5865__B1 _2486_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_943 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8527__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6409__A2 mod.Data_Mem.F_M.MRAM\[12\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_497 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8572__D _0076_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7209__I1 mod.Data_Mem.F_M.MRAM\[2\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_1101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_1123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_1156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6968__I0 _3405_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5985__S _1515_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6042__B1 _2656_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2180 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4800_ _1464_ _1466_ _1469_ _1470_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XTAP_2191 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5780_ _2403_ _2404_ _2405_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4731_ _1347_ _1385_ _1401_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_147_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7450_ _3698_ _0433_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6345__A1 _1608_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4662_ mod.Arithmetic.CN.I_in\[38\] _1332_ _1251_ _1333_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_163_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6401_ _2418_ mod.Data_Mem.F_M.MRAM\[780\]\[0\] _3010_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_7381_ mod.Data_Mem.F_M.MRAM\[773\]\[7\] _3664_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_134_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4593_ _0786_ _0855_ _0628_ _1265_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__8057__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6332_ _2868_ _2935_ _2943_ _2944_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_127_193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_116_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6499__I2 mod.Data_Mem.F_M.MRAM\[781\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6263_ _1737_ _2876_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_103_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7504__I _3321_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8002_ _0211_ net1 mod.Data_Mem.F_M.MRAM\[13\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5214_ _1790_ _1879_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_88_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6194_ _2765_ _2807_ _2808_ _2809_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_57_604 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5145_ _1503_ _1811_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_96_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5024__I _1579_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5608__B1 _2243_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5076_ mod.Data_Mem.F_M.MRAM\[17\]\[2\] mod.Data_Mem.F_M.MRAM\[16\]\[2\] _1519_ _1743_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_84_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4027_ _0638_ mod.Arithmetic.I_out\[72\] _0703_ _0704_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_72_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_1201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_1212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7620__I1 mod.Data_Mem.F_M.MRAM\[787\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5978_ _2385_ mod.Data_Mem.F_M.MRAM\[782\]\[5\] _2597_ _2598_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_7717_ _3852_ _0546_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4929_ _1597_ _1598_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_7648_ mod.Data_Mem.F_M.MRAM\[790\]\[0\] _3818_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_20_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__6336__A1 _2846_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_20_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7579_ _3777_ _0483_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_101_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7615__S _3798_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_1216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3942__I _0619_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_169_1126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_16_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_43_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_157_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_129_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6590__A4 _3179_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6327__A1 _2904_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6327__B2 _2267_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_145_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_11_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5925__I1 _1901_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5550__A2 mod.Data_Mem.F_M.MRAM\[30\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7827__A1 _3908_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8567__D _0071_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_504 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7917__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_526 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6350__I1 _1996_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_548 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_604 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_59_90 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_1193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_773 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5066__A1 mod.Data_Mem.F_M.MRAM\[6\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4683__I mod.Arithmetic.CN.I_in\[53\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_787 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6950_ _3235_ _3407_ _3374_ _3408_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_82_938 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_75_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5901_ mod.Data_Mem.F_M.MRAM\[18\]\[3\] mod.Data_Mem.F_M.MRAM\[19\]\[3\] _2522_ _2523_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_6881_ mod.Data_Mem.F_M.MRAM\[4\]\[0\] _3363_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_35_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_62_640 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5832_ _2447_ _2455_ _2456_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_62_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6566__A1 _1966_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8551_ _0055_ net1 mod.Data_Mem.F_M.out_data\[31\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_72_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_868 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5763_ _2101_ _2388_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_124_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7502_ _3729_ mod.Data_Mem.F_M.MRAM\[781\]\[6\] _3726_ _3730_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4714_ _1349_ _1384_ _1385_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__6318__A1 _2886_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8482_ _0578_ net1 mod.Data_Mem.F_M.MRAM\[798\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5694_ _2280_ _2140_ _2320_ _2322_ _2323_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
X_7433_ mod.Data_Mem.F_M.MRAM\[777\]\[1\] _3690_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4645_ _1061_ _1313_ _1315_ _1316_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_135_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_7364_ _3655_ _0390_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_162_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4576_ _1241_ _1247_ _1248_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_6315_ _2872_ _1958_ _2927_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_115_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7295_ _3555_ _3606_ _3614_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_89_526 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_859 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6246_ _2858_ _2221_ _1664_ _2859_ _2860_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_130_166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_924 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6177_ _2199_ _2682_ _2792_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_97_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5910__C _1800_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5128_ _1530_ _1795_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_85_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2905 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5059_ _1698_ _1723_ _1726_ _1727_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_2916 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_426 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2927 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_84_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2938 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2949 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_168_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6006__B1 _2624_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4280__A2 _0646_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_504 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6557__A1 _2312_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8222__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3937__I _0614_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5080__I1 mod.Data_Mem.F_M.MRAM\[18\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_166_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5780__A2 _2404_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4969__S _1636_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8372__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5907__I1 mod.Data_Mem.F_M.MRAM\[17\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7345__S _3643_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5532__A2 _2172_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_1160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_1019 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_84 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_122_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_430 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5296__A1 _1622_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_110_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5820__C _2443_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_90_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4008__I _0638_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_1126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_44_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6548__A1 _1491_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_1137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_1197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_12_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_31 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4430_ _1089_ _1102_ _1103_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_144_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4361_ _0781_ _0854_ _0856_ _1033_ _1034_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_113_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6100_ _2710_ _2689_ _2716_ _2717_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_7080_ mod.Data_Mem.F_M.MRAM\[21\]\[3\] _3487_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__7520__I0 _3645_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4292_ _0870_ _0878_ _0879_ _0966_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or3_1
XFILLER_115_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6893__I mod.Data_Mem.F_M.MRAM\[4\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6031_ _2506_ mod.Data_Mem.F_M.MRAM\[788\]\[7\] _2648_ _2649_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_98_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_356 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_367 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_7982_ mod.Instr_Mem.instruction\[7\] net2 net1 mod.P1.instr_reg\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XANTENNA__5302__I _1965_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_584 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8245__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5834__I0 mod.Data_Mem.F_M.MRAM\[30\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6933_ _3396_ _0218_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_70_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_35_651 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_29 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_74_1204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6864_ _3354_ _0191_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6539__A1 _2522_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7587__I0 _3782_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_168_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_50_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5815_ _2422_ _2439_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__8395__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6795_ _3299_ _3313_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_50_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8534_ _0038_ net1 mod.Data_Mem.F_M.out_data\[46\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_148_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5746_ _2362_ _2364_ _2365_ _2355_ _2370_ _2371_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_22_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5762__A2 mod.Data_Mem.F_M.MRAM\[768\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7339__I0 _3531_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8465_ _0561_ net1 mod.Data_Mem.F_M.MRAM\[796\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5677_ _2135_ mod.Data_Mem.F_M.MRAM\[797\]\[3\] _2307_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_124_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7416_ _3681_ _0416_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_11_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4628_ _1185_ _1093_ _1184_ _1299_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_8396_ _0492_ net1 mod.Data_Mem.F_M.MRAM\[786\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__5514__A2 mod.Data_Mem.F_M.MRAM\[798\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_163_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7347_ _3618_ mod.Data_Mem.F_M.MRAM\[771\]\[6\] _3643_ _3647_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4559_ _1227_ _1230_ _1231_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_89_312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7278_ _3601_ _0358_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__7511__I0 _3638_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_6229_ _2838_ _2842_ _2843_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_890 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_765 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_85_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_724 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5212__I _1580_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2702 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2713 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2724 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2735 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2746 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5450__A1 _2097_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2757 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2768 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2779 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_610 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_13_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5368__B _1863_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5738__C1 _2361_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_41_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5087__C _1616_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_1061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_167_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_1083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__4961__B1 _1624_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_1078 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_5_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5505__A2 mod.Data_Mem.F_M.MRAM\[30\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7750__I0 _3749_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8118__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput4 net4 io_out[17] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XFILLER_134_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_150_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7502__I0 _3729_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_987 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8268__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_62_1152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_49_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4492__A2 _1076_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_1196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_787 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5441__A1 _2080_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_1002 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5600_ mod.Data_Mem.F_M.MRAM\[797\]\[4\] _2221_ _1749_ mod.Data_Mem.F_M.MRAM\[796\]\[4\]
+ _2236_ _2237_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XFILLER_34_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6580_ mod.I_addr\[4\] _3178_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5744__A2 _2368_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_157_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5531_ _2170_ mod.Data_Mem.F_M.MRAM\[798\]\[0\] mod.Data_Mem.F_M.MRAM\[799\]\[0\]
+ _2171_ _2172_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_75_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_8_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8250_ _0346_ net1 mod.Data_Mem.F_M.MRAM\[31\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5462_ _2108_ _2110_ _2111_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__5347__I2 mod.Data_Mem.F_M.MRAM\[789\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_145_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7201_ _3508_ mod.Data_Mem.F_M.MRAM\[29\]\[5\] _3553_ _3558_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4413_ _1002_ _1022_ _1086_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_8181_ _0291_ net1 mod.Data_Mem.F_M.MRAM\[3\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_114_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5393_ _2048_ _2054_ _1775_ _2055_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_7132_ _3452_ mod.Data_Mem.F_M.MRAM\[19\]\[2\] _3513_ _3516_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_119_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4344_ _1017_ _1018_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_67_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_1085 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6457__B1 _2642_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_59_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7063_ _3478_ _0266_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_98_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4275_ _0866_ _0886_ _0949_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_115_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6556__C _2108_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6014_ _2512_ mod.Data_Mem.F_M.MRAM\[21\]\[6\] _2633_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5680__A1 _2306_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_584 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5032__I _1562_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2009 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_94_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7965_ _0191_ net1 mod.Data_Mem.F_M.MRAM\[779\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_36_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_43_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5967__I _2214_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1319 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_78_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6916_ _3256_ mod.Data_Mem.F_M.MRAM\[13\]\[6\] _3381_ _3384_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_7896_ _0122_ net1 mod.Data_Mem.F_M.MRAM\[27\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__5983__A2 _1934_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_23_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_643 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6847_ _3259_ mod.Data_Mem.F_M.MRAM\[769\]\[7\] _3336_ _3346_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_51_985 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_149_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6778_ _3299_ _3300_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__6783__I1 _3303_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6798__I net8 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8517_ net185 net1 mod.Data_Mem.F_M.out_data\[61\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5729_ _1812_ _1553_ _2354_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_136_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_109_759 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8448_ _0544_ net1 mod.Data_Mem.F_M.MRAM\[794\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_108_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5499__A1 _1879_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_8379_ _0475_ net1 mod.Data_Mem.F_M.MRAM\[784\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_117_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4171__A1 _0665_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8410__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_1174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_751 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6299__I0 _2232_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_968 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3200 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8560__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3211 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3222 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_3233 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7799__I0 _3322_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3244 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_133_96 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2510 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3255 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2521 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2532 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_716 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5877__I _2395_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5423__A1 _2080_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2543 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2554 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2565 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1820 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_749 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1831 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2576 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5974__A2 _2590_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2587 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1842 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2598 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1853 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3985__A1 _0650_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1864 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1875 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_1886 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1897 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6501__I _2203_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_155_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_10_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6151__A2 _1649_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8090__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4162__A1 _0635_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4956__I _1489_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_151_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_151_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4060_ mod.Arithmetic.CN.I_in\[14\] _0737_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_110_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5662__A1 _2168_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_1061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_83_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_830 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_149_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_52_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4217__A2 mod.Arithmetic.CN.I_in\[34\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4962_ _1630_ _0000_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_7750_ _3749_ mod.Data_Mem.F_M.MRAM\[796\]\[2\] _3867_ _3870_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__5965__A2 _2143_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_248 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6701_ _3249_ mod.Data_Mem.F_M.MRAM\[28\]\[4\] _3250_ _3251_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_51_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7681_ _3834_ _0528_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4893_ _1561_ _1562_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_20_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6632_ _3206_ _0107_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_20_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6563_ mod.Data_Mem.F_M.MRAM\[780\]\[7\] _1674_ _3107_ _3164_ _2698_ _3165_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_118_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4640__B _1061_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5228__S _1892_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5514_ _2138_ mod.Data_Mem.F_M.MRAM\[798\]\[7\] _2155_ _2156_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_8302_ _0398_ net1 mod.Data_Mem.F_M.MRAM\[773\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__6411__I _2376_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8433__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6494_ _3096_ _3097_ _3098_ _3099_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_8233_ _0329_ net1 mod.Data_Mem.F_M.MRAM\[2\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5445_ _2078_ _2093_ _2094_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5027__I _1571_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4153__A1 _0828_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8164_ mod.Data_Mem.F_M.out_data\[74\] net2 net1 mod.Arithmetic.I_out\[74\] vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_5376_ _2023_ _2030_ _2031_ _2037_ _1899_ _2038_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
X_7115_ _3505_ _0291_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__8583__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_160_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6059__S _2295_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4327_ _0993_ _0999_ _1001_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_141_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_8095_ mod.Data_Mem.F_M.out_data\[5\] net2 net1 mod.Arithmetic.ACTI.x\[5\] vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_86_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5328__S1 _1882_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6286__C _1866_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_646 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7046_ _3452_ mod.Data_Mem.F_M.MRAM\[1\]\[2\] _3469_ _3470_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_75_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4258_ _0929_ _0931_ _0932_ _0933_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_101_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_86_167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5653__A1 _2280_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4189_ _0819_ _0851_ _0864_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_27_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_167_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4208__A2 _0814_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5405__A1 _1724_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_103_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1116 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_70_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1127 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_7948_ _0174_ net1 mod.Data_Mem.F_M.MRAM\[789\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1149 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3967__A1 _0643_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_169_924 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7879_ _0105_ net1 mod.Data_Mem.F_M.MRAM\[26\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_51_771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7618__S _3801_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_793 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_169_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_168_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5708__A2 mod.Data_Mem.F_M.MRAM\[29\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__3945__I _0622_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4042__S _0702_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4392__A1 _1061_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4392__B2 _0871_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6133__A2 _2747_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5892__A1 _2511_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7950__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5644__A1 _2275_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6692__I0 _3243_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6991__I _3234_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_830 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_690 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3030 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3041 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_19_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_3052 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3063 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8306__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3074 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3085 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2340 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3096 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2351 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_535 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2362 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2373 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2384 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1051 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1650 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2395 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1661 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1672 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7528__S _3745_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1683 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1694 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8456__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_1049 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4383__A1 _0634_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5275__C _1563_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_154_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7263__S _3590_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5230_ mod.Data_Mem.F_M.MRAM\[17\]\[4\] mod.Data_Mem.F_M.MRAM\[16\]\[4\] _1894_ _1895_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__4135__A1 _0644_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_1180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5883__A1 _2423_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_5161_ mod.Data_Mem.F_M.MRAM\[785\]\[3\] mod.Data_Mem.F_M.MRAM\[784\]\[3\] _1685_
+ _1827_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_69_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4112_ _0743_ _0778_ _0788_ _0789_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_68_145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_765 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5092_ _1597_ _1759_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_84_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_56_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4043_ _0710_ _0712_ _0719_ _0630_ _0720_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_84_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_830 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_690 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_37_532 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_513 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7802_ _3899_ _0584_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_80_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5994_ _2587_ mod.Data_Mem.F_M.MRAM\[788\]\[6\] _2612_ _2613_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_64_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6060__A1 _2565_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_169_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7733_ _3860_ _0554_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_36_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4945_ _1561_ _1614_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_75_1162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4610__A2 _1257_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6342__S _1738_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7664_ mod.Data_Mem.F_M.MRAM\[791\]\[0\] _3826_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4876_ mod.Data_Mem.F_M.MRAM\[3\]\[0\] _1539_ _1531_ _1544_ _1545_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_60_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5246__S0 _1910_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6615_ mod.Data_Mem.F_M.MRAM\[24\]\[3\] _3198_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_7595_ _3788_ _0488_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_119_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6546_ _3049_ _2341_ _2500_ _2615_ _2616_ _2568_ _3149_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_146_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6477_ _2189_ _3083_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__7163__I1 mod.Data_Mem.F_M.MRAM\[12\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7973__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5428_ _2083_ _0017_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_8216_ _0317_ net1 mod.Data_Mem.F_M.MRAM\[22\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5359_ _2000_ _2021_ _2022_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_8147_ mod.Data_Mem.F_M.out_data\[57\] net2 net1 mod.Arithmetic.CN.I_in\[57\] vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_99_270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_134_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_99_292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8078_ mod.P3.Res\[6\] net2 net1 net9 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_82_1188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_988 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_21 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8329__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5477__I1 mod.Data_Mem.F_M.MRAM\[31\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7029_ _3458_ _0252_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_75_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_800 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_43_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8479__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_749 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_31 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_169_765 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6354__A2 mod.Data_Mem.F_M.MRAM\[15\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_7_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_7_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_165_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4117__A1 _0673_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_879 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_79_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_79_911 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5865__A1 _2449_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4668__A2 _1338_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_124_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_105_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_966 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_540 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8099__RN net2 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5617__A1 _1737_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5331__S _1708_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_11 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_77 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6968__I1 mod.Data_Mem.F_M.MRAM\[15\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6042__A1 _2423_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_1168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6042__B2 _2464_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2170 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2181 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2192 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4730_ _1349_ _1400_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_1480 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1491 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4661_ _1090_ _1330_ _1331_ _1332_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_159_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6345__A2 _1989_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6400_ _2499_ _3009_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4356__A1 _0775_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7996__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7380_ _3663_ _0398_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5553__B1 _2159_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_156_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4592_ _0786_ _0799_ _0857_ _1263_ _1264_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_70_1092 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6331_ _2867_ _2942_ _2943_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_157_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_155_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6262_ _1655_ _1880_ _2875_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__6499__I3 _1901_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5856__A1 _2281_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8001_ _0210_ net1 mod.Data_Mem.F_M.MRAM\[13\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5213_ mod.Data_Mem.F_M.MRAM\[1\]\[4\] mod.Data_Mem.F_M.MRAM\[0\]\[4\] _1877_ _1878_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_88_229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6193_ _2180_ _1735_ _2808_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_69_432 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_752 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5144_ mod.Data_Mem.F_M.MRAM\[6\]\[3\] _1645_ _1808_ _1809_ _1557_ _1810_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_69_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5608__A1 _2225_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5608__B2 _2177_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5075_ _1524_ _1742_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_56_126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_852 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6281__A1 _2886_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4026_ _0702_ _0703_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__6136__I _1564_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6033__A1 _2097_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6584__A2 _3179_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5977_ _1933_ mod.Data_Mem.F_M.MRAM\[783\]\[5\] _2597_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_40_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7716_ mod.Data_Mem.F_M.MRAM\[794\]\[2\] _3852_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_100_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4928_ _1594_ _1596_ _1597_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_165_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7647_ _3817_ _0511_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4859_ _1521_ _1492_ _1528_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__8001__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7578_ _3765_ mod.Data_Mem.F_M.MRAM\[785\]\[3\] _3773_ _3777_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_147_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6529_ _2534_ _3123_ _3132_ _0077_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__7836__A2 mod.I_addr\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8151__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5847__A1 _2358_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_1050 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_678 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_48_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5151__S _1816_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_169_1116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_169_1149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7869__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_1021 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_169_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6327__A2 mod.Data_Mem.F_M.MRAM\[783\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4338__A1 _0914_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_125_610 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5326__S _1609_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7827__A2 _3913_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_153_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_112_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_113_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_505 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_538 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_538 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_1161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_120_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5066__A2 _1601_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5310__I0 mod.Data_Mem.F_M.MRAM\[3\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_980 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5900_ _1609_ _2522_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_93_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6880_ _3362_ _0199_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6015__A1 _2548_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5831_ _2449_ _2450_ _2451_ _2357_ _2453_ _2454_ _2455_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_61_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8024__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_1121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8550_ _0054_ net1 mod.Data_Mem.F_M.out_data\[30\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5762_ _2385_ mod.Data_Mem.F_M.MRAM\[768\]\[0\] _2386_ _2387_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_7501_ _3318_ _3729_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_72_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4713_ _1363_ _1383_ _1384_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_147_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5693_ _2321_ mod.Data_Mem.F_M.MRAM\[796\]\[4\] _2311_ _2322_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_8481_ _0577_ net1 mod.Data_Mem.F_M.MRAM\[798\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_33_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_163_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7432_ _3689_ _0424_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4644_ _1063_ _1178_ _1314_ _1315_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__5526__B1 _2159_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8174__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7363_ mod.Data_Mem.F_M.MRAM\[772\]\[6\] _3655_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4575_ _1242_ _1246_ _1247_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_128_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5129__I0 _1781_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6314_ _2924_ _2925_ _2926_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_7294_ _1770_ _3609_ _3613_ _0362_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_116_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_157_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6245_ _2129_ mod.Data_Mem.F_M.MRAM\[783\]\[3\] mod.Data_Mem.F_M.MRAM\[782\]\[3\]
+ _2070_ _2859_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_44_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4501__A1 _0678_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6176_ _2749_ _2758_ _2791_ _2374_ _0065_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_69_251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5127_ _1791_ mod.Data_Mem.F_M.MRAM\[785\]\[2\] _1793_ _1794_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__4874__I _1542_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_969 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5058_ _1725_ _1726_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_2906 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2917 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2928 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4009_ _0684_ mod.Arithmetic.I_out\[73\] mod.Arithmetic.I_out\[72\] _0685_ _0686_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XTAP_2939 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_1032 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_169_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7054__I0 _3460_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6006__B2 _2611_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4280__A3 _0809_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6557__A2 _2508_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4542__C _0980_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8517__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7626__S _3801_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_166_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_153_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_107_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3953__I mod.Arithmetic.CN.I_in\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_49_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_1014 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4740__A1 _1407_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_84_1069 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6493__A1 _2345_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5296__A2 _1959_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_914 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_497 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_48_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_102_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6245__A1 _2129_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6245__B2 _2070_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_788 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_213 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__8047__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_1121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_1116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_1149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4559__A1 _1227_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5220__A2 _1883_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8197__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7536__S _3745_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_145_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5508__B1 _2150_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__8578__D _0594_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4031__I0 _0682_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_1201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5374__I3 _2035_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_1212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4360_ _0780_ _0795_ _1033_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_141_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4291_ _0953_ _0955_ _0964_ _0965_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XANTENNA__7520__I1 mod.Data_Mem.F_M.MRAM\[782\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6030_ _2428_ mod.Data_Mem.F_M.MRAM\[789\]\[7\] _2648_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__6484__A1 _3030_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_819 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_66_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7981_ _0207_ net1 mod.Data_Mem.F_M.MRAM\[4\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__5834__I1 _1632_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_82_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6932_ _3395_ mod.Data_Mem.F_M.MRAM\[14\]\[2\] _3391_ _3396_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_35_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_19 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__7036__I0 _3462_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_1216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6863_ mod.Data_Mem.F_M.MRAM\[779\]\[7\] _3354_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_62_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6539__A2 mod.Data_Mem.F_M.MRAM\[781\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5814_ mod.Data_Mem.F_M.MRAM\[782\]\[1\] mod.Data_Mem.F_M.MRAM\[783\]\[1\] _1918_
+ _2438_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_34_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6794_ _3311_ _3312_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_37_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8533_ _0037_ net1 mod.Data_Mem.F_M.out_data\[45\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5745_ _2366_ _2369_ _2370_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_50_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7339__I1 mod.Data_Mem.F_M.MRAM\[771\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6350__S _1713_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8464_ _0560_ net1 mod.Data_Mem.F_M.MRAM\[796\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__4970__A1 _1635_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5676_ _2132_ _2306_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_135_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_148_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_108_429 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7415_ mod.Data_Mem.F_M.MRAM\[776\]\[0\] _3681_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4869__I _1537_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4627_ _1185_ _1093_ _1184_ _1298_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_8395_ _0491_ net1 mod.Data_Mem.F_M.MRAM\[786\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_7346_ _3646_ _0381_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4558_ _1228_ _1229_ _1230_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_117_985 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7277_ mod.Data_Mem.F_M.MRAM\[5\]\[6\] _3601_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4489_ _1048_ _1077_ _1161_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_104_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6475__A1 _3004_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6228_ mod.Data_Mem.F_M.MRAM\[13\]\[3\] _1729_ _2840_ _2841_ _2842_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_44_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_1042 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_880 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6159_ _2713_ _2775_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_66_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_97_390 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_891 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4537__C _0983_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_79_1127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_980 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_57_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_58_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2703 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2714 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4109__I mod.Arithmetic.ACTI.x\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2725 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2736 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2747 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2758 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2769 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7907__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_158_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_1051 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_51_1013 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_1193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_90_1073 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4961__A1 _1491_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_716 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4961__B2 _1629_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_108_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_123_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput5 net5 io_out[18] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XFILLER_123_933 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7502__I1 mod.Data_Mem.F_M.MRAM\[781\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6466__A1 _3063_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_1164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5403__I _1501_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6218__A1 _2212_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_48_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7018__I0 _3450_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5441__A2 _2077_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_972 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_674 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_1014 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_290 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_9_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5530_ _1782_ _2171_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_117_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5461_ _2109_ _2110_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_68_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_7200_ _3557_ _0324_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4412_ _1002_ _1022_ _1085_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__4704__A1 _0641_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8180_ _0290_ net1 mod.Data_Mem.F_M.MRAM\[3\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5392_ _2012_ _2051_ _2053_ _1822_ _2054_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_160_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_158_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7131_ _3515_ _0297_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_114_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4343_ mod.Arithmetic.CN.I_in\[59\] _1017_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_113_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4180__A2 mod.P2.Rout_reg\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8212__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6457__A1 mod.Data_Mem.F_M.MRAM\[13\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7062_ mod.Data_Mem.F_M.MRAM\[20\]\[2\] _3478_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_67_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6457__B2 mod.Data_Mem.F_M.MRAM\[1\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_465 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4274_ _0946_ _0947_ _0948_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_99_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6013_ _2549_ mod.Data_Mem.F_M.MRAM\[20\]\[6\] _2632_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_67_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6209__A1 _2186_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7257__I0 mod.Data_Mem.F_M.MRAM\[31\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5680__A2 _2309_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8362__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7964_ _0190_ net1 mod.Data_Mem.F_M.MRAM\[779\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__7009__I0 _3405_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1309 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_78_1160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6915_ _3383_ _0213_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_35_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_739 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7895_ _0121_ net1 mod.Data_Mem.F_M.MRAM\[27\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_35_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_168_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6846_ _3345_ _0182_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__3994__A2 _0670_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4092__C _0768_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5196__A1 _1552_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_167_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6777_ _3294_ _3296_ _3298_ _3299_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_22_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3989_ _0663_ _0665_ _0666_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_8516_ net186 net1 mod.Data_Mem.F_M.out_data\[60\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_10_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5728_ _2352_ _2353_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_164_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8447_ _0543_ net1 mod.Data_Mem.F_M.MRAM\[793\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5659_ _1914_ _2290_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_108_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5499__A2 mod.Data_Mem.F_M.MRAM\[30\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_163_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5743__I0 mod.Data_Mem.F_M.MRAM\[2\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8378_ _0474_ net1 mod.Data_Mem.F_M.MRAM\[784\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_105_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7329_ _3272_ _3296_ _3634_ _3635_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_105_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_1006 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6448__A1 _3004_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6299__I1 _2237_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7248__I0 mod.Data_Mem.F_M.MRAM\[31\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3201 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3212 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3223 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7799__I1 mod.Data_Mem.F_M.MRAM\[798\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3234 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_533 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3245 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2500 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3256 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2511 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2522 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2533 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5423__A2 _2077_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2544 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2555 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1810 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2566 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1821 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2577 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1832 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2588 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1843 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1854 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2599 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3985__A2 _0661_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1865 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_1119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1876 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_159_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1887 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5187__A1 _1845_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1898 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_105_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_41_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6384__B1 mod.Data_Mem.F_M.MRAM\[14\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5982__I0 mod.Data_Mem.F_M.MRAM\[770\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_154_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_127_535 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6003__B _2621_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8235__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5734__I0 mod.Data_Mem.F_M.MRAM\[14\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_1204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4162__A2 mod.Arithmetic.CN.I_in\[49\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5334__S _1894_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7487__I0 _3718_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__8385__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5133__I _1799_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5662__A2 _2292_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4972__I _1639_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_64_588 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4961_ _1491_ _1498_ _1560_ _1624_ _1629_ _1630_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai32_1
XANTENNA__5965__A3 _2145_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6700_ _3236_ _3250_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_32_430 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7680_ mod.Data_Mem.F_M.MRAM\[792\]\[0\] _3834_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA_output4_I net4 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4892_ _1554_ _1504_ _1561_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_60_761 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6631_ mod.Data_Mem.F_M.MRAM\[26\]\[3\] _3206_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_149_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6562_ _2385_ mod.Data_Mem.F_M.MRAM\[768\]\[7\] _3164_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_146_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_1085 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8301_ _0397_ net1 mod.Data_Mem.F_M.MRAM\[773\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5513_ _1715_ mod.Data_Mem.F_M.MRAM\[799\]\[7\] _2155_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_6493_ _2345_ mod.Data_Mem.F_M.MRAM\[2\]\[4\] _2440_ _2569_ _3098_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_145_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8232_ _0328_ net1 mod.Data_Mem.F_M.MRAM\[2\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_133_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5444_ _2092_ _1619_ _2093_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_69_1159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_161_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4153__A2 _0820_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8163_ mod.Data_Mem.F_M.out_data\[73\] net2 net1 mod.Arithmetic.I_out\[73\] vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_5375_ _1888_ _2036_ _1621_ _2037_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__5244__S _1908_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7114_ _3454_ mod.Data_Mem.F_M.MRAM\[3\]\[3\] _3501_ _3505_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__7478__I0 _3645_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_603 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4326_ _0993_ _0999_ _1000_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_8094_ mod.Data_Mem.F_M.out_data\[4\] net2 net1 mod.Arithmetic.ACTI.x\[4\] vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_102_936 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7045_ _3465_ _3469_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_4257_ _0824_ _0929_ _0931_ _0932_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_101_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5653__A2 _2121_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_714 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_67_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_68_894 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4188_ _0821_ _0822_ _0669_ _0850_ _0863_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_132_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_67_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_28_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_67_393 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5199__B _1625_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1106 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1117 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_7947_ _0173_ net1 mod.Data_Mem.F_M.MRAM\[789\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__8108__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1128 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5956__A3 _2576_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1139 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_24_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_430 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3967__A2 mod.Arithmetic.CN.I_in\[16\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7878_ _0104_ net1 mod.Data_Mem.F_M.MRAM\[26\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_169_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_6829_ _3334_ _3335_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_51_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8258__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_31 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_10_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4392__A2 _1063_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_31 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3961__I mod.Arithmetic.CN.I_in\[16\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_151_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_105_752 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_120_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6692__I1 mod.Data_Mem.F_M.MRAM\[28\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_319 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_500 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6493__B _2440_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_3020 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3031 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3042 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3053 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3064 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3075 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2330 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3086 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2341 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2352 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_3097 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2363 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2374 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2385 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1640 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2396 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1651 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1662 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1673 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1684 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6357__B1 mod.Data_Mem.F_M.MRAM\[782\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1695 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_800 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_155_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5580__A1 _2061_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5128__I _1530_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7544__S _3752_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4032__I mod.Arithmetic.CN.I_in\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5064__S _1636_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_603 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5160_ _1663_ _1826_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_68_1192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5883__A2 _2131_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_123_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_1056 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4111_ _0740_ _0766_ _0788_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_96_433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_97_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5091_ _1757_ mod.Data_Mem.F_M.MRAM\[31\]\[2\] _1721_ mod.Data_Mem.F_M.MRAM\[15\]\[2\]
+ _1758_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_110_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4042_ _0685_ _0718_ _0702_ _0719_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_68_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_639 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7801_ mod.Data_Mem.F_M.MRAM\[7\]\[0\] _3899_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_80_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_37_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_536 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5993_ _2588_ mod.Data_Mem.F_M.MRAM\[789\]\[6\] _2612_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_52_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_91_193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7732_ mod.Data_Mem.F_M.MRAM\[795\]\[2\] _3860_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_52_569 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4944_ mod.Data_Mem.F_M.MRAM\[785\]\[0\] mod.Data_Mem.F_M.MRAM\[784\]\[0\] _1612_
+ _1613_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_75_1152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8400__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_75_1185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7663_ _3825_ _0519_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4875_ mod.Data_Mem.F_M.MRAM\[6\]\[0\] _1540_ _1543_ _1544_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_60_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5239__S _1903_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_162_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6899__A1 mod.Data_Mem.F_M.dest\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6422__I _2429_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6614_ _3197_ _0098_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5246__S1 _1805_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7594_ _3771_ mod.Data_Mem.F_M.MRAM\[786\]\[0\] _3787_ _3788_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_137_129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_118_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6545_ _2611_ _2627_ _3144_ _2211_ _3147_ _3148_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XANTENNA__8550__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4374__A2 _0974_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_888 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6476_ _2184_ _3079_ _3081_ _3082_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_8215_ _0316_ net1 mod.Data_Mem.F_M.MRAM\[22\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__4126__A2 _0648_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5323__A1 mod.Data_Mem.F_M.MRAM\[15\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5427_ _1802_ _2082_ _2083_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_133_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_47_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8146_ mod.Data_Mem.F_M.out_data\[56\] net2 net1 mod.Arithmetic.CN.I_in\[56\] vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_99_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_160_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5358_ _2001_ _2007_ _2020_ _1927_ _1629_ _2021_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_88_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_1167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4309_ _0650_ mod.Arithmetic.CN.I_in\[43\] _0983_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_102_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8077_ mod.P3.Res\[5\] net2 net1 net8 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_5289_ _1579_ _1953_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_101_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_788 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_33 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_500 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7028_ _3456_ mod.Data_Mem.F_M.MRAM\[18\]\[4\] _3457_ _3458_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_74_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_87_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_28_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6051__A2 _2668_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8080__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_169_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3956__I _0632_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_168_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_51_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_169_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_128_118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4988__S _1519_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_11_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_836 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_139_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_155_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5865__A2 _2485_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_891 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_639 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_820 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5411__I _2069_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8423__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_1114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_62_823 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7539__S _3752_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2160 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6042__A2 _2655_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2171 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_81 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2182 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_62_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2193 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_21_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_61_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1470 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8573__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1481 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1492 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4660_ _0651_ mod.Arithmetic.CN.I_in\[35\] _1090_ _1330_ _1331_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XANTENNA__5553__A1 _2169_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4591_ _0785_ _0795_ _1263_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5553__B2 _2192_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6330_ _2240_ _2243_ _2938_ _2941_ _1964_ _2759_ _2942_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_116_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_116_858 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6261_ _2872_ _1876_ _2873_ _2874_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_89_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8000_ _0209_ net1 mod.Data_Mem.F_M.MRAM\[13\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5212_ _1580_ _1877_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_88_219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5856__A2 mod.Data_Mem.F_M.MRAM\[772\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6192_ _1742_ _1739_ _2807_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_97_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_123_390 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5143_ _1543_ _1809_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_69_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_904 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7801__I mod.Data_Mem.F_M.MRAM\[7\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_85_915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5608__A2 _2240_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5074_ _1732_ _1733_ _1736_ _1740_ _1741_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_56_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_4025_ mod.Arithmetic.CN.I_in\[23\] _0677_ _0694_ _0700_ _0701_ _0702_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_4
XANTENNA__6417__I _2092_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_801 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7605__I0 _3754_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_25_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_71_119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6033__A2 mod.Data_Mem.F_M.MRAM\[786\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5976_ _2381_ _2596_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_7715_ _3851_ _0545_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_52_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_539 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4927_ _1595_ _1494_ _1596_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_7646_ mod.Data_Mem.F_M.MRAM\[788\]\[7\] _3817_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__7940__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4858_ _1526_ _1527_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_21_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_166_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_119_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7577_ _3776_ _0482_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4789_ _1329_ _1345_ _1458_ _1459_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_165_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6528_ _2626_ _3129_ _3131_ _2079_ _3132_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_107_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_162_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_109_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6459_ _2619_ mod.Data_Mem.F_M.MRAM\[0\]\[2\] _3066_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_106_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_161_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8129_ mod.Data_Mem.F_M.out_data\[39\] net2 net1 mod.Arithmetic.CN.I_in\[39\] vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_130_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__8446__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_1087 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_21_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_169_1128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4283__A1 _0875_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_44_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_1033 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5783__A1 _2406_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_169_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_165_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4310__I _0983_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_3_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_539 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_390 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_81 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6438__S _2512_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5342__S _1908_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_959 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_94_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5310__I1 mod.Data_Mem.F_M.MRAM\[2\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5830_ _2354_ _2454_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_61_130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_962 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7963__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7763__A2 _3705_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6566__A3 _3167_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_995 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_1111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5761_ _1954_ mod.Data_Mem.F_M.MRAM\[769\]\[0\] _2386_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__5774__A1 _2398_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_7500_ _3728_ _0453_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_124_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4712_ _1365_ _1382_ _1383_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_72_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8480_ _0576_ net1 mod.Data_Mem.F_M.MRAM\[798\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5692_ _1593_ _2321_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_148_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6318__A3 _2929_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_1188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7431_ mod.Data_Mem.F_M.MRAM\[777\]\[0\] _3689_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__8319__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4643_ mod.Arithmetic.CN.I_in\[30\] _1314_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5526__A1 _2081_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5526__B2 _2165_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_147_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6700__I _3236_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7362_ _3654_ _0389_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_128_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4574_ _1243_ _1245_ _1246_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_144_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6313_ _1826_ _1952_ _2873_ _2925_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__5129__I1 _1786_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7293_ _3612_ _3606_ _3613_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_118_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__8469__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6244_ mod.Data_Mem.F_M.MRAM\[781\]\[3\] _2858_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__5385__S0 _1829_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4501__A2 mod.Arithmetic.CN.I_in\[20\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6175_ _1670_ _2778_ _2784_ _2790_ _2743_ _2791_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XFILLER_97_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5126_ _1715_ _1792_ _1793_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_85_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_745 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6147__I _2713_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5057_ _1724_ _1725_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_2907 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2918 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4008_ _0638_ _0685_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XANTENNA__4804__A3 _1473_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2929 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6006__A2 _2622_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7054__I1 mod.Data_Mem.F_M.MRAM\[1\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_1055 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_13_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4017__A1 _0679_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_675 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_984 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6557__A3 _2668_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_1200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_40_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5959_ _2457_ _2578_ _1536_ _2362_ _2579_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XANTENNA__5000__B _1622_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7994__RN net2 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7629_ _2013_ _3804_ _3808_ _0502_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_5_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_147_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_31 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_1004 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_1184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_106_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_432 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8171__RN net2 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6493__A2 mod.Data_Mem.F_M.MRAM\[2\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_75_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6245__A2 mod.Data_Mem.F_M.MRAM\[783\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_929 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4256__A1 _0621_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7986__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_1133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_962 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_984 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_1019 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4559__A2 _1230_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_169_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7985__RN net2 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5508__A1 _2119_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5508__B2 _2133_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6181__A1 _2687_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4031__I1 mod.Arithmetic.I_out\[74\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_430 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5136__I _1695_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_153_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_99_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4290_ _0962_ _0963_ _0964_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_125_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5367__S0 _1881_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5580__B _2217_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8594__D _0610_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6484__A2 _2514_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8162__RN net2 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5072__S _1647_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_358 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_67_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_121_680 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_7980_ _0206_ net1 mod.Data_Mem.F_M.MRAM\[4\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_94_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5295__I0 _1950_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6931_ _3242_ _3395_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5995__A1 _2214_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4798__A2 _1176_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7036__I1 mod.Data_Mem.F_M.MRAM\[18\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6862_ _3353_ _0190_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_35_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_781 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5813_ _2321_ _1709_ _2436_ _2437_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_90_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_161_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8141__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5747__A1 _2353_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6793_ net7 _3311_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_22_358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8532_ _0036_ net1 mod.Data_Mem.F_M.out_data\[44\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5744_ _2367_ _2368_ _2369_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_124_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_8463_ _0559_ net1 mod.Data_Mem.F_M.MRAM\[795\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5675_ _2076_ _2304_ _2166_ _2305_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__4970__A2 _1637_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8291__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7414_ _3680_ _0415_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_129_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4626_ _1293_ _1296_ _1297_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__6172__A1 _1734_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8394_ _0490_ net1 mod.Data_Mem.F_M.MRAM\[786\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_159_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_151_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7345_ _3645_ mod.Data_Mem.F_M.MRAM\[771\]\[5\] _3643_ _3646_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_132_901 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5046__I _1578_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4557_ mod.Arithmetic.CN.I_in\[53\] _1114_ _1116_ _1229_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_116_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7276_ _3600_ _0357_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4488_ _1048_ _1077_ _1160_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__4885__I mod.Data_Mem.F_M.src\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8153__RN net2 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6475__A2 _3080_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6227_ _1619_ _2702_ _2841_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_106_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6158_ _2761_ _1665_ _2774_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6227__A2 _2702_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5109_ mod.Data_Mem.F_M.MRAM\[783\]\[2\] _1775_ _1776_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_73_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6089_ _1494_ _1542_ _2706_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_100_875 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2704 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2715 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2726 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2737 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2748 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2759 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_25_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5738__A1 _2112_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_41_645 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_678 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5665__B _2259_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4961__A2 _1498_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3964__I _0640_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_739 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_5_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_166_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_430 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput6 net6 io_out[19] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XFILLER_135_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8144__RN net2 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8014__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_163_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_49_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6218__A2 _2219_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5977__A1 _1933_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8164__CLK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5729__A1 _1812_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_20_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_34_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_180 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_191 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_158_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6154__A1 _1751_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5460_ _2069_ _2064_ _2109_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_133_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4411_ _0988_ _1083_ _1084_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__4704__A2 mod.Arithmetic.ACTI.x\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5391_ _1704_ _2052_ _2053_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_99_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_1032 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7130_ _3450_ mod.Data_Mem.F_M.MRAM\[19\]\[1\] _3513_ _3515_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4342_ _1007_ _1015_ _1016_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_154_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_67_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6457__A2 _2382_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7061_ _3477_ _0265_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__8135__RN net2 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6701__I0 _3249_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4273_ _0866_ _0886_ _0947_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_6012_ mod.Data_Mem.F_M.MRAM\[16\]\[6\] mod.Data_Mem.F_M.MRAM\[17\]\[6\] _2418_ _2631_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_100_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
.ends

