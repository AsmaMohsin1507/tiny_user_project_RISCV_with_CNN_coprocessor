magic
tech gf180mcuC
magscale 1 5
timestamp 1670001947
<< obsm1 >>
rect 672 855 69328 68529
<< metal2 >>
rect 672 69600 728 69900
rect 1344 69600 1400 69900
rect 2016 69600 2072 69900
rect 2688 69600 2744 69900
rect 3360 69600 3416 69900
rect 4032 69600 4088 69900
rect 4704 69600 4760 69900
rect 5376 69600 5432 69900
rect 6048 69600 6104 69900
rect 6720 69600 6776 69900
rect 7392 69600 7448 69900
rect 8064 69600 8120 69900
rect 8736 69600 8792 69900
rect 9408 69600 9464 69900
rect 10080 69600 10136 69900
rect 10752 69600 10808 69900
rect 11424 69600 11480 69900
rect 12096 69600 12152 69900
rect 12768 69600 12824 69900
rect 13440 69600 13496 69900
rect 14112 69600 14168 69900
rect 14784 69600 14840 69900
rect 15456 69600 15512 69900
rect 16128 69600 16184 69900
rect 16800 69600 16856 69900
rect 17472 69600 17528 69900
rect 18144 69600 18200 69900
rect 18816 69600 18872 69900
rect 19488 69600 19544 69900
rect 20160 69600 20216 69900
rect 20832 69600 20888 69900
rect 21504 69600 21560 69900
rect 22176 69600 22232 69900
rect 22848 69600 22904 69900
rect 23520 69600 23576 69900
rect 24192 69600 24248 69900
rect 24864 69600 24920 69900
rect 25536 69600 25592 69900
rect 26208 69600 26264 69900
rect 26880 69600 26936 69900
rect 27552 69600 27608 69900
rect 28224 69600 28280 69900
rect 28896 69600 28952 69900
rect 29568 69600 29624 69900
rect 30240 69600 30296 69900
rect 30912 69600 30968 69900
rect 31584 69600 31640 69900
rect 32256 69600 32312 69900
rect 32928 69600 32984 69900
rect 33600 69600 33656 69900
rect 34272 69600 34328 69900
rect 34944 69600 35000 69900
rect 35616 69600 35672 69900
rect 36288 69600 36344 69900
rect 36960 69600 37016 69900
rect 37632 69600 37688 69900
rect 38304 69600 38360 69900
rect 38976 69600 39032 69900
rect 39648 69600 39704 69900
rect 40320 69600 40376 69900
rect 40992 69600 41048 69900
rect 41664 69600 41720 69900
rect 42336 69600 42392 69900
rect 43008 69600 43064 69900
rect 43680 69600 43736 69900
rect 44352 69600 44408 69900
rect 45024 69600 45080 69900
rect 45696 69600 45752 69900
rect 46368 69600 46424 69900
rect 47040 69600 47096 69900
rect 47712 69600 47768 69900
rect 48384 69600 48440 69900
rect 49056 69600 49112 69900
rect 49728 69600 49784 69900
rect 50400 69600 50456 69900
rect 51072 69600 51128 69900
rect 51744 69600 51800 69900
rect 52416 69600 52472 69900
rect 53088 69600 53144 69900
rect 53760 69600 53816 69900
rect 54432 69600 54488 69900
rect 55104 69600 55160 69900
rect 55776 69600 55832 69900
rect 56448 69600 56504 69900
rect 57120 69600 57176 69900
rect 57792 69600 57848 69900
rect 58464 69600 58520 69900
rect 59136 69600 59192 69900
rect 59808 69600 59864 69900
rect 60480 69600 60536 69900
rect 61152 69600 61208 69900
rect 61824 69600 61880 69900
rect 62496 69600 62552 69900
rect 63168 69600 63224 69900
rect 63840 69600 63896 69900
rect 64512 69600 64568 69900
rect 65184 69600 65240 69900
rect 65856 69600 65912 69900
rect 66528 69600 66584 69900
rect 67200 69600 67256 69900
rect 67872 69600 67928 69900
rect 68544 69600 68600 69900
rect 69216 69600 69272 69900
rect 69888 69600 69944 69900
rect 0 100 56 400
rect 672 100 728 400
rect 1344 100 1400 400
rect 2016 100 2072 400
rect 2688 100 2744 400
rect 3360 100 3416 400
rect 4032 100 4088 400
rect 4704 100 4760 400
rect 5376 100 5432 400
rect 6048 100 6104 400
rect 6720 100 6776 400
rect 7392 100 7448 400
rect 8064 100 8120 400
rect 8736 100 8792 400
rect 9408 100 9464 400
rect 10080 100 10136 400
rect 10752 100 10808 400
rect 11424 100 11480 400
rect 12096 100 12152 400
rect 12768 100 12824 400
rect 13440 100 13496 400
rect 14112 100 14168 400
rect 14784 100 14840 400
rect 15456 100 15512 400
rect 16128 100 16184 400
rect 16800 100 16856 400
rect 17472 100 17528 400
rect 18144 100 18200 400
rect 18816 100 18872 400
rect 19488 100 19544 400
rect 20160 100 20216 400
rect 20832 100 20888 400
rect 21504 100 21560 400
rect 22176 100 22232 400
rect 22848 100 22904 400
rect 23520 100 23576 400
rect 24192 100 24248 400
rect 24864 100 24920 400
rect 25536 100 25592 400
rect 26208 100 26264 400
rect 26880 100 26936 400
rect 27552 100 27608 400
rect 28224 100 28280 400
rect 28896 100 28952 400
rect 29568 100 29624 400
rect 30240 100 30296 400
rect 30912 100 30968 400
rect 31584 100 31640 400
rect 32256 100 32312 400
rect 32928 100 32984 400
rect 33600 100 33656 400
rect 34272 100 34328 400
rect 34944 100 35000 400
rect 35616 100 35672 400
rect 36288 100 36344 400
rect 36960 100 37016 400
rect 37632 100 37688 400
rect 38304 100 38360 400
rect 38976 100 39032 400
rect 39648 100 39704 400
rect 40320 100 40376 400
rect 40992 100 41048 400
rect 41664 100 41720 400
rect 42336 100 42392 400
rect 43008 100 43064 400
rect 43680 100 43736 400
rect 44352 100 44408 400
rect 45024 100 45080 400
rect 45696 100 45752 400
rect 46368 100 46424 400
rect 47040 100 47096 400
rect 47712 100 47768 400
rect 48384 100 48440 400
rect 49056 100 49112 400
rect 49728 100 49784 400
rect 50400 100 50456 400
rect 51072 100 51128 400
rect 51744 100 51800 400
rect 52416 100 52472 400
rect 53088 100 53144 400
rect 53760 100 53816 400
rect 54432 100 54488 400
rect 55104 100 55160 400
rect 55776 100 55832 400
rect 56448 100 56504 400
rect 57120 100 57176 400
rect 57792 100 57848 400
rect 58464 100 58520 400
rect 59136 100 59192 400
rect 59808 100 59864 400
rect 60480 100 60536 400
rect 61152 100 61208 400
rect 61824 100 61880 400
rect 62496 100 62552 400
rect 63168 100 63224 400
rect 63840 100 63896 400
rect 64512 100 64568 400
rect 65184 100 65240 400
rect 65856 100 65912 400
rect 66528 100 66584 400
rect 67200 100 67256 400
rect 67872 100 67928 400
rect 68544 100 68600 400
rect 69216 100 69272 400
<< obsm2 >>
rect 14 69930 69538 69935
rect 14 69570 642 69930
rect 758 69570 1314 69930
rect 1430 69570 1986 69930
rect 2102 69570 2658 69930
rect 2774 69570 3330 69930
rect 3446 69570 4002 69930
rect 4118 69570 4674 69930
rect 4790 69570 5346 69930
rect 5462 69570 6018 69930
rect 6134 69570 6690 69930
rect 6806 69570 7362 69930
rect 7478 69570 8034 69930
rect 8150 69570 8706 69930
rect 8822 69570 9378 69930
rect 9494 69570 10050 69930
rect 10166 69570 10722 69930
rect 10838 69570 11394 69930
rect 11510 69570 12066 69930
rect 12182 69570 12738 69930
rect 12854 69570 13410 69930
rect 13526 69570 14082 69930
rect 14198 69570 14754 69930
rect 14870 69570 15426 69930
rect 15542 69570 16098 69930
rect 16214 69570 16770 69930
rect 16886 69570 17442 69930
rect 17558 69570 18114 69930
rect 18230 69570 18786 69930
rect 18902 69570 19458 69930
rect 19574 69570 20130 69930
rect 20246 69570 20802 69930
rect 20918 69570 21474 69930
rect 21590 69570 22146 69930
rect 22262 69570 22818 69930
rect 22934 69570 23490 69930
rect 23606 69570 24162 69930
rect 24278 69570 24834 69930
rect 24950 69570 25506 69930
rect 25622 69570 26178 69930
rect 26294 69570 26850 69930
rect 26966 69570 27522 69930
rect 27638 69570 28194 69930
rect 28310 69570 28866 69930
rect 28982 69570 29538 69930
rect 29654 69570 30210 69930
rect 30326 69570 30882 69930
rect 30998 69570 31554 69930
rect 31670 69570 32226 69930
rect 32342 69570 32898 69930
rect 33014 69570 33570 69930
rect 33686 69570 34242 69930
rect 34358 69570 34914 69930
rect 35030 69570 35586 69930
rect 35702 69570 36258 69930
rect 36374 69570 36930 69930
rect 37046 69570 37602 69930
rect 37718 69570 38274 69930
rect 38390 69570 38946 69930
rect 39062 69570 39618 69930
rect 39734 69570 40290 69930
rect 40406 69570 40962 69930
rect 41078 69570 41634 69930
rect 41750 69570 42306 69930
rect 42422 69570 42978 69930
rect 43094 69570 43650 69930
rect 43766 69570 44322 69930
rect 44438 69570 44994 69930
rect 45110 69570 45666 69930
rect 45782 69570 46338 69930
rect 46454 69570 47010 69930
rect 47126 69570 47682 69930
rect 47798 69570 48354 69930
rect 48470 69570 49026 69930
rect 49142 69570 49698 69930
rect 49814 69570 50370 69930
rect 50486 69570 51042 69930
rect 51158 69570 51714 69930
rect 51830 69570 52386 69930
rect 52502 69570 53058 69930
rect 53174 69570 53730 69930
rect 53846 69570 54402 69930
rect 54518 69570 55074 69930
rect 55190 69570 55746 69930
rect 55862 69570 56418 69930
rect 56534 69570 57090 69930
rect 57206 69570 57762 69930
rect 57878 69570 58434 69930
rect 58550 69570 59106 69930
rect 59222 69570 59778 69930
rect 59894 69570 60450 69930
rect 60566 69570 61122 69930
rect 61238 69570 61794 69930
rect 61910 69570 62466 69930
rect 62582 69570 63138 69930
rect 63254 69570 63810 69930
rect 63926 69570 64482 69930
rect 64598 69570 65154 69930
rect 65270 69570 65826 69930
rect 65942 69570 66498 69930
rect 66614 69570 67170 69930
rect 67286 69570 67842 69930
rect 67958 69570 68514 69930
rect 68630 69570 69186 69930
rect 69302 69570 69538 69930
rect 14 430 69538 69570
rect 86 400 642 430
rect 758 400 1314 430
rect 1430 400 1986 430
rect 2102 400 2658 430
rect 2774 400 3330 430
rect 3446 400 4002 430
rect 4118 400 4674 430
rect 4790 400 5346 430
rect 5462 400 6018 430
rect 6134 400 6690 430
rect 6806 400 7362 430
rect 7478 400 8034 430
rect 8150 400 8706 430
rect 8822 400 9378 430
rect 9494 400 10050 430
rect 10166 400 10722 430
rect 10838 400 11394 430
rect 11510 400 12066 430
rect 12182 400 12738 430
rect 12854 400 13410 430
rect 13526 400 14082 430
rect 14198 400 14754 430
rect 14870 400 15426 430
rect 15542 400 16098 430
rect 16214 400 16770 430
rect 16886 400 17442 430
rect 17558 400 18114 430
rect 18230 400 18786 430
rect 18902 400 19458 430
rect 19574 400 20130 430
rect 20246 400 20802 430
rect 20918 400 21474 430
rect 21590 400 22146 430
rect 22262 400 22818 430
rect 22934 400 23490 430
rect 23606 400 24162 430
rect 24278 400 24834 430
rect 24950 400 25506 430
rect 25622 400 26178 430
rect 26294 400 26850 430
rect 26966 400 27522 430
rect 27638 400 28194 430
rect 28310 400 28866 430
rect 28982 400 29538 430
rect 29654 400 30210 430
rect 30326 400 30882 430
rect 30998 400 31554 430
rect 31670 400 32226 430
rect 32342 400 32898 430
rect 33014 400 33570 430
rect 33686 400 34242 430
rect 34358 400 34914 430
rect 35030 400 35586 430
rect 35702 400 36258 430
rect 36374 400 36930 430
rect 37046 400 37602 430
rect 37718 400 38274 430
rect 38390 400 38946 430
rect 39062 400 39618 430
rect 39734 400 40290 430
rect 40406 400 40962 430
rect 41078 400 41634 430
rect 41750 400 42306 430
rect 42422 400 42978 430
rect 43094 400 43650 430
rect 43766 400 44322 430
rect 44438 400 44994 430
rect 45110 400 45666 430
rect 45782 400 46338 430
rect 46454 400 47010 430
rect 47126 400 47682 430
rect 47798 400 48354 430
rect 48470 400 49026 430
rect 49142 400 49698 430
rect 49814 400 50370 430
rect 50486 400 51042 430
rect 51158 400 51714 430
rect 51830 400 52386 430
rect 52502 400 53058 430
rect 53174 400 53730 430
rect 53846 400 54402 430
rect 54518 400 55074 430
rect 55190 400 55746 430
rect 55862 400 56418 430
rect 56534 400 57090 430
rect 57206 400 57762 430
rect 57878 400 58434 430
rect 58550 400 59106 430
rect 59222 400 59778 430
rect 59894 400 60450 430
rect 60566 400 61122 430
rect 61238 400 61794 430
rect 61910 400 62466 430
rect 62582 400 63138 430
rect 63254 400 63810 430
rect 63926 400 64482 430
rect 64598 400 65154 430
rect 65270 400 65826 430
rect 65942 400 66498 430
rect 66614 400 67170 430
rect 67286 400 67842 430
rect 67958 400 68514 430
rect 68630 400 69186 430
rect 69302 400 69538 430
<< metal3 >>
rect 100 69888 400 69944
rect 100 69216 400 69272
rect 69600 69216 69900 69272
rect 100 68544 400 68600
rect 69600 68544 69900 68600
rect 100 67872 400 67928
rect 69600 67872 69900 67928
rect 100 67200 400 67256
rect 69600 67200 69900 67256
rect 100 66528 400 66584
rect 69600 66528 69900 66584
rect 100 65856 400 65912
rect 69600 65856 69900 65912
rect 100 65184 400 65240
rect 69600 65184 69900 65240
rect 100 64512 400 64568
rect 69600 64512 69900 64568
rect 100 63840 400 63896
rect 69600 63840 69900 63896
rect 100 63168 400 63224
rect 69600 63168 69900 63224
rect 100 62496 400 62552
rect 69600 62496 69900 62552
rect 100 61824 400 61880
rect 69600 61824 69900 61880
rect 100 61152 400 61208
rect 69600 61152 69900 61208
rect 100 60480 400 60536
rect 69600 60480 69900 60536
rect 100 59808 400 59864
rect 69600 59808 69900 59864
rect 100 59136 400 59192
rect 69600 59136 69900 59192
rect 100 58464 400 58520
rect 69600 58464 69900 58520
rect 100 57792 400 57848
rect 69600 57792 69900 57848
rect 100 57120 400 57176
rect 69600 57120 69900 57176
rect 100 56448 400 56504
rect 69600 56448 69900 56504
rect 100 55776 400 55832
rect 69600 55776 69900 55832
rect 100 55104 400 55160
rect 69600 55104 69900 55160
rect 100 54432 400 54488
rect 69600 54432 69900 54488
rect 100 53760 400 53816
rect 69600 53760 69900 53816
rect 100 53088 400 53144
rect 69600 53088 69900 53144
rect 100 52416 400 52472
rect 69600 52416 69900 52472
rect 100 51744 400 51800
rect 69600 51744 69900 51800
rect 100 51072 400 51128
rect 69600 51072 69900 51128
rect 100 50400 400 50456
rect 69600 50400 69900 50456
rect 100 49728 400 49784
rect 69600 49728 69900 49784
rect 100 49056 400 49112
rect 69600 49056 69900 49112
rect 100 48384 400 48440
rect 69600 48384 69900 48440
rect 100 47712 400 47768
rect 69600 47712 69900 47768
rect 100 47040 400 47096
rect 69600 47040 69900 47096
rect 100 46368 400 46424
rect 69600 46368 69900 46424
rect 100 45696 400 45752
rect 69600 45696 69900 45752
rect 100 45024 400 45080
rect 69600 45024 69900 45080
rect 100 44352 400 44408
rect 69600 44352 69900 44408
rect 100 43680 400 43736
rect 69600 43680 69900 43736
rect 100 43008 400 43064
rect 69600 43008 69900 43064
rect 100 42336 400 42392
rect 69600 42336 69900 42392
rect 100 41664 400 41720
rect 69600 41664 69900 41720
rect 100 40992 400 41048
rect 69600 40992 69900 41048
rect 100 40320 400 40376
rect 69600 40320 69900 40376
rect 100 39648 400 39704
rect 69600 39648 69900 39704
rect 100 38976 400 39032
rect 69600 38976 69900 39032
rect 100 38304 400 38360
rect 69600 38304 69900 38360
rect 100 37632 400 37688
rect 69600 37632 69900 37688
rect 100 36960 400 37016
rect 69600 36960 69900 37016
rect 100 36288 400 36344
rect 69600 36288 69900 36344
rect 100 35616 400 35672
rect 69600 35616 69900 35672
rect 100 34944 400 35000
rect 69600 34944 69900 35000
rect 100 34272 400 34328
rect 69600 34272 69900 34328
rect 100 33600 400 33656
rect 69600 33600 69900 33656
rect 100 32928 400 32984
rect 69600 32928 69900 32984
rect 100 32256 400 32312
rect 69600 32256 69900 32312
rect 100 31584 400 31640
rect 69600 31584 69900 31640
rect 100 30912 400 30968
rect 69600 30912 69900 30968
rect 100 30240 400 30296
rect 69600 30240 69900 30296
rect 100 29568 400 29624
rect 69600 29568 69900 29624
rect 100 28896 400 28952
rect 69600 28896 69900 28952
rect 100 28224 400 28280
rect 69600 28224 69900 28280
rect 100 27552 400 27608
rect 69600 27552 69900 27608
rect 100 26880 400 26936
rect 69600 26880 69900 26936
rect 100 26208 400 26264
rect 69600 26208 69900 26264
rect 100 25536 400 25592
rect 69600 25536 69900 25592
rect 100 24864 400 24920
rect 69600 24864 69900 24920
rect 100 24192 400 24248
rect 69600 24192 69900 24248
rect 100 23520 400 23576
rect 69600 23520 69900 23576
rect 100 22848 400 22904
rect 69600 22848 69900 22904
rect 100 22176 400 22232
rect 69600 22176 69900 22232
rect 100 21504 400 21560
rect 69600 21504 69900 21560
rect 100 20832 400 20888
rect 69600 20832 69900 20888
rect 100 20160 400 20216
rect 69600 20160 69900 20216
rect 100 19488 400 19544
rect 69600 19488 69900 19544
rect 100 18816 400 18872
rect 69600 18816 69900 18872
rect 100 18144 400 18200
rect 69600 18144 69900 18200
rect 100 17472 400 17528
rect 69600 17472 69900 17528
rect 100 16800 400 16856
rect 69600 16800 69900 16856
rect 100 16128 400 16184
rect 69600 16128 69900 16184
rect 100 15456 400 15512
rect 69600 15456 69900 15512
rect 100 14784 400 14840
rect 69600 14784 69900 14840
rect 100 14112 400 14168
rect 69600 14112 69900 14168
rect 100 13440 400 13496
rect 69600 13440 69900 13496
rect 100 12768 400 12824
rect 69600 12768 69900 12824
rect 100 12096 400 12152
rect 69600 12096 69900 12152
rect 100 11424 400 11480
rect 69600 11424 69900 11480
rect 100 10752 400 10808
rect 69600 10752 69900 10808
rect 100 10080 400 10136
rect 69600 10080 69900 10136
rect 100 9408 400 9464
rect 69600 9408 69900 9464
rect 100 8736 400 8792
rect 69600 8736 69900 8792
rect 100 8064 400 8120
rect 69600 8064 69900 8120
rect 100 7392 400 7448
rect 69600 7392 69900 7448
rect 100 6720 400 6776
rect 69600 6720 69900 6776
rect 100 6048 400 6104
rect 69600 6048 69900 6104
rect 100 5376 400 5432
rect 69600 5376 69900 5432
rect 100 4704 400 4760
rect 69600 4704 69900 4760
rect 100 4032 400 4088
rect 69600 4032 69900 4088
rect 100 3360 400 3416
rect 69600 3360 69900 3416
rect 100 2688 400 2744
rect 69600 2688 69900 2744
rect 100 2016 400 2072
rect 69600 2016 69900 2072
rect 100 1344 400 1400
rect 69600 1344 69900 1400
rect 100 672 400 728
rect 69600 672 69900 728
rect 69600 0 69900 56
<< obsm3 >>
rect 9 69858 70 69930
rect 430 69858 69650 69930
rect 9 69302 69650 69858
rect 9 69186 70 69302
rect 430 69186 69570 69302
rect 9 68630 69650 69186
rect 9 68514 70 68630
rect 430 68514 69570 68630
rect 9 67958 69650 68514
rect 9 67842 70 67958
rect 430 67842 69570 67958
rect 9 67286 69650 67842
rect 9 67170 70 67286
rect 430 67170 69570 67286
rect 9 66614 69650 67170
rect 9 66498 70 66614
rect 430 66498 69570 66614
rect 9 65942 69650 66498
rect 9 65826 70 65942
rect 430 65826 69570 65942
rect 9 65270 69650 65826
rect 9 65154 70 65270
rect 430 65154 69570 65270
rect 9 64598 69650 65154
rect 9 64482 70 64598
rect 430 64482 69570 64598
rect 9 63926 69650 64482
rect 9 63810 70 63926
rect 430 63810 69570 63926
rect 9 63254 69650 63810
rect 9 63138 70 63254
rect 430 63138 69570 63254
rect 9 62582 69650 63138
rect 9 62466 70 62582
rect 430 62466 69570 62582
rect 9 61910 69650 62466
rect 9 61794 70 61910
rect 430 61794 69570 61910
rect 9 61238 69650 61794
rect 9 61122 70 61238
rect 430 61122 69570 61238
rect 9 60566 69650 61122
rect 9 60450 70 60566
rect 430 60450 69570 60566
rect 9 59894 69650 60450
rect 9 59778 70 59894
rect 430 59778 69570 59894
rect 9 59222 69650 59778
rect 9 59106 70 59222
rect 430 59106 69570 59222
rect 9 58550 69650 59106
rect 9 58434 70 58550
rect 430 58434 69570 58550
rect 9 57878 69650 58434
rect 9 57762 70 57878
rect 430 57762 69570 57878
rect 9 57206 69650 57762
rect 9 57090 70 57206
rect 430 57090 69570 57206
rect 9 56534 69650 57090
rect 9 56418 70 56534
rect 430 56418 69570 56534
rect 9 55862 69650 56418
rect 9 55746 70 55862
rect 430 55746 69570 55862
rect 9 55190 69650 55746
rect 9 55074 70 55190
rect 430 55074 69570 55190
rect 9 54518 69650 55074
rect 9 54402 70 54518
rect 430 54402 69570 54518
rect 9 53846 69650 54402
rect 9 53730 70 53846
rect 430 53730 69570 53846
rect 9 53174 69650 53730
rect 9 53058 70 53174
rect 430 53058 69570 53174
rect 9 52502 69650 53058
rect 9 52386 70 52502
rect 430 52386 69570 52502
rect 9 51830 69650 52386
rect 9 51714 70 51830
rect 430 51714 69570 51830
rect 9 51158 69650 51714
rect 9 51042 70 51158
rect 430 51042 69570 51158
rect 9 50486 69650 51042
rect 9 50370 70 50486
rect 430 50370 69570 50486
rect 9 49814 69650 50370
rect 9 49698 70 49814
rect 430 49698 69570 49814
rect 9 49142 69650 49698
rect 9 49026 70 49142
rect 430 49026 69570 49142
rect 9 48470 69650 49026
rect 9 48354 70 48470
rect 430 48354 69570 48470
rect 9 47798 69650 48354
rect 9 47682 70 47798
rect 430 47682 69570 47798
rect 9 47126 69650 47682
rect 9 47010 70 47126
rect 430 47010 69570 47126
rect 9 46454 69650 47010
rect 9 46338 70 46454
rect 430 46338 69570 46454
rect 9 45782 69650 46338
rect 9 45666 70 45782
rect 430 45666 69570 45782
rect 9 45110 69650 45666
rect 9 44994 70 45110
rect 430 44994 69570 45110
rect 9 44438 69650 44994
rect 9 44322 70 44438
rect 430 44322 69570 44438
rect 9 43766 69650 44322
rect 9 43650 70 43766
rect 430 43650 69570 43766
rect 9 43094 69650 43650
rect 9 42978 70 43094
rect 430 42978 69570 43094
rect 9 42422 69650 42978
rect 9 42306 70 42422
rect 430 42306 69570 42422
rect 9 41750 69650 42306
rect 9 41634 70 41750
rect 430 41634 69570 41750
rect 9 41078 69650 41634
rect 9 40962 70 41078
rect 430 40962 69570 41078
rect 9 40406 69650 40962
rect 9 40290 70 40406
rect 430 40290 69570 40406
rect 9 39734 69650 40290
rect 9 39618 70 39734
rect 430 39618 69570 39734
rect 9 39062 69650 39618
rect 9 38946 70 39062
rect 430 38946 69570 39062
rect 9 38390 69650 38946
rect 9 38274 70 38390
rect 430 38274 69570 38390
rect 9 37718 69650 38274
rect 9 37602 70 37718
rect 430 37602 69570 37718
rect 9 37046 69650 37602
rect 9 36930 70 37046
rect 430 36930 69570 37046
rect 9 36374 69650 36930
rect 9 36258 70 36374
rect 430 36258 69570 36374
rect 9 35702 69650 36258
rect 9 35586 70 35702
rect 430 35586 69570 35702
rect 9 35030 69650 35586
rect 9 34914 70 35030
rect 430 34914 69570 35030
rect 9 34358 69650 34914
rect 9 34242 70 34358
rect 430 34242 69570 34358
rect 9 33686 69650 34242
rect 9 33570 70 33686
rect 430 33570 69570 33686
rect 9 33014 69650 33570
rect 9 32898 70 33014
rect 430 32898 69570 33014
rect 9 32342 69650 32898
rect 9 32226 70 32342
rect 430 32226 69570 32342
rect 9 31670 69650 32226
rect 9 31554 70 31670
rect 430 31554 69570 31670
rect 9 30998 69650 31554
rect 9 30882 70 30998
rect 430 30882 69570 30998
rect 9 30326 69650 30882
rect 9 30210 70 30326
rect 430 30210 69570 30326
rect 9 29654 69650 30210
rect 9 29538 70 29654
rect 430 29538 69570 29654
rect 9 28982 69650 29538
rect 9 28866 70 28982
rect 430 28866 69570 28982
rect 9 28310 69650 28866
rect 9 28194 70 28310
rect 430 28194 69570 28310
rect 9 27638 69650 28194
rect 9 27522 70 27638
rect 430 27522 69570 27638
rect 9 26966 69650 27522
rect 9 26850 70 26966
rect 430 26850 69570 26966
rect 9 26294 69650 26850
rect 9 26178 70 26294
rect 430 26178 69570 26294
rect 9 25622 69650 26178
rect 9 25506 70 25622
rect 430 25506 69570 25622
rect 9 24950 69650 25506
rect 9 24834 70 24950
rect 430 24834 69570 24950
rect 9 24278 69650 24834
rect 9 24162 70 24278
rect 430 24162 69570 24278
rect 9 23606 69650 24162
rect 9 23490 70 23606
rect 430 23490 69570 23606
rect 9 22934 69650 23490
rect 9 22818 70 22934
rect 430 22818 69570 22934
rect 9 22262 69650 22818
rect 9 22146 70 22262
rect 430 22146 69570 22262
rect 9 21590 69650 22146
rect 9 21474 70 21590
rect 430 21474 69570 21590
rect 9 20918 69650 21474
rect 9 20802 70 20918
rect 430 20802 69570 20918
rect 9 20246 69650 20802
rect 9 20130 70 20246
rect 430 20130 69570 20246
rect 9 19574 69650 20130
rect 9 19458 70 19574
rect 430 19458 69570 19574
rect 9 18902 69650 19458
rect 9 18786 70 18902
rect 430 18786 69570 18902
rect 9 18230 69650 18786
rect 9 18114 70 18230
rect 430 18114 69570 18230
rect 9 17558 69650 18114
rect 9 17442 70 17558
rect 430 17442 69570 17558
rect 9 16886 69650 17442
rect 9 16770 70 16886
rect 430 16770 69570 16886
rect 9 16214 69650 16770
rect 9 16098 70 16214
rect 430 16098 69570 16214
rect 9 15542 69650 16098
rect 9 15426 70 15542
rect 430 15426 69570 15542
rect 9 14870 69650 15426
rect 9 14754 70 14870
rect 430 14754 69570 14870
rect 9 14198 69650 14754
rect 9 14082 70 14198
rect 430 14082 69570 14198
rect 9 13526 69650 14082
rect 9 13410 70 13526
rect 430 13410 69570 13526
rect 9 12854 69650 13410
rect 9 12738 70 12854
rect 430 12738 69570 12854
rect 9 12182 69650 12738
rect 9 12066 70 12182
rect 430 12066 69570 12182
rect 9 11510 69650 12066
rect 9 11394 70 11510
rect 430 11394 69570 11510
rect 9 10838 69650 11394
rect 9 10722 70 10838
rect 430 10722 69570 10838
rect 9 10166 69650 10722
rect 9 10050 70 10166
rect 430 10050 69570 10166
rect 9 9494 69650 10050
rect 9 9378 70 9494
rect 430 9378 69570 9494
rect 9 8822 69650 9378
rect 9 8706 70 8822
rect 430 8706 69570 8822
rect 9 8150 69650 8706
rect 9 8034 70 8150
rect 430 8034 69570 8150
rect 9 7478 69650 8034
rect 9 7362 70 7478
rect 430 7362 69570 7478
rect 9 6806 69650 7362
rect 9 6690 70 6806
rect 430 6690 69570 6806
rect 9 6134 69650 6690
rect 9 6018 70 6134
rect 430 6018 69570 6134
rect 9 5462 69650 6018
rect 9 5346 70 5462
rect 430 5346 69570 5462
rect 9 4790 69650 5346
rect 9 4674 70 4790
rect 430 4674 69570 4790
rect 9 4118 69650 4674
rect 9 4002 70 4118
rect 430 4002 69570 4118
rect 9 3446 69650 4002
rect 9 3330 70 3446
rect 430 3330 69570 3446
rect 9 2774 69650 3330
rect 9 2658 70 2774
rect 430 2658 69570 2774
rect 9 2102 69650 2658
rect 9 1986 70 2102
rect 430 1986 69570 2102
rect 9 1430 69650 1986
rect 9 1314 70 1430
rect 430 1314 69570 1430
rect 9 758 69650 1314
rect 9 642 70 758
rect 430 642 69570 758
rect 9 518 69650 642
<< metal4 >>
rect 2224 1538 2384 68238
rect 9904 1538 10064 68238
rect 17584 1538 17744 68238
rect 25264 1538 25424 68238
rect 32944 1538 33104 68238
rect 40624 1538 40784 68238
rect 48304 1538 48464 68238
rect 55984 1538 56144 68238
rect 63664 1538 63824 68238
<< obsm4 >>
rect 10990 1508 17554 58287
rect 17774 1508 25234 58287
rect 25454 1508 32914 58287
rect 33134 1508 40594 58287
rect 40814 1508 48274 58287
rect 48494 1508 55954 58287
rect 56174 1508 63634 58287
rect 63854 1508 68754 58287
rect 10990 513 68754 1508
<< labels >>
rlabel metal3 s 100 48384 400 48440 6 io_in[0]
port 1 nsew signal input
rlabel metal3 s 100 49056 400 49112 6 io_in[10]
port 2 nsew signal input
rlabel metal3 s 100 24192 400 24248 6 io_in[11]
port 3 nsew signal input
rlabel metal3 s 100 42336 400 42392 6 io_in[12]
port 4 nsew signal input
rlabel metal3 s 100 28896 400 28952 6 io_in[13]
port 5 nsew signal input
rlabel metal3 s 100 24864 400 24920 6 io_in[14]
port 6 nsew signal input
rlabel metal2 s 36960 69600 37016 69900 6 io_in[15]
port 7 nsew signal input
rlabel metal3 s 69600 14112 69900 14168 6 io_in[16]
port 8 nsew signal input
rlabel metal3 s 69600 65856 69900 65912 6 io_in[17]
port 9 nsew signal input
rlabel metal2 s 47040 69600 47096 69900 6 io_in[18]
port 10 nsew signal input
rlabel metal2 s 68544 100 68600 400 6 io_in[19]
port 11 nsew signal input
rlabel metal2 s 8736 69600 8792 69900 6 io_in[1]
port 12 nsew signal input
rlabel metal2 s 55776 69600 55832 69900 6 io_in[20]
port 13 nsew signal input
rlabel metal2 s 49056 100 49112 400 6 io_in[21]
port 14 nsew signal input
rlabel metal2 s 69888 69600 69944 69900 6 io_in[22]
port 15 nsew signal input
rlabel metal3 s 69600 60480 69900 60536 6 io_in[23]
port 16 nsew signal input
rlabel metal2 s 57792 100 57848 400 6 io_in[24]
port 17 nsew signal input
rlabel metal2 s 9408 100 9464 400 6 io_in[25]
port 18 nsew signal input
rlabel metal3 s 100 58464 400 58520 6 io_in[26]
port 19 nsew signal input
rlabel metal3 s 100 47712 400 47768 6 io_in[27]
port 20 nsew signal input
rlabel metal3 s 100 54432 400 54488 6 io_in[28]
port 21 nsew signal input
rlabel metal3 s 100 43680 400 43736 6 io_in[29]
port 22 nsew signal input
rlabel metal3 s 69600 69216 69900 69272 6 io_in[2]
port 23 nsew signal input
rlabel metal2 s 45696 100 45752 400 6 io_in[30]
port 24 nsew signal input
rlabel metal3 s 100 29568 400 29624 6 io_in[31]
port 25 nsew signal input
rlabel metal2 s 59136 100 59192 400 6 io_in[32]
port 26 nsew signal input
rlabel metal3 s 100 7392 400 7448 6 io_in[33]
port 27 nsew signal input
rlabel metal3 s 100 62496 400 62552 6 io_in[34]
port 28 nsew signal input
rlabel metal2 s 62496 69600 62552 69900 6 io_in[35]
port 29 nsew signal input
rlabel metal3 s 69600 61824 69900 61880 6 io_in[36]
port 30 nsew signal input
rlabel metal3 s 69600 53088 69900 53144 6 io_in[37]
port 31 nsew signal input
rlabel metal3 s 69600 68544 69900 68600 6 io_in[3]
port 32 nsew signal input
rlabel metal3 s 69600 31584 69900 31640 6 io_in[4]
port 33 nsew signal input
rlabel metal3 s 100 13440 400 13496 6 io_in[5]
port 34 nsew signal input
rlabel metal3 s 69600 13440 69900 13496 6 io_in[6]
port 35 nsew signal input
rlabel metal2 s 57120 69600 57176 69900 6 io_in[7]
port 36 nsew signal input
rlabel metal3 s 100 32256 400 32312 6 io_in[8]
port 37 nsew signal input
rlabel metal3 s 100 36288 400 36344 6 io_in[9]
port 38 nsew signal input
rlabel metal3 s 69600 49056 69900 49112 6 io_oeb[0]
port 39 nsew signal output
rlabel metal3 s 69600 45024 69900 45080 6 io_oeb[10]
port 40 nsew signal output
rlabel metal2 s 2688 69600 2744 69900 6 io_oeb[11]
port 41 nsew signal output
rlabel metal2 s 43008 100 43064 400 6 io_oeb[12]
port 42 nsew signal output
rlabel metal3 s 100 18144 400 18200 6 io_oeb[13]
port 43 nsew signal output
rlabel metal2 s 63840 100 63896 400 6 io_oeb[14]
port 44 nsew signal output
rlabel metal2 s 44352 69600 44408 69900 6 io_oeb[15]
port 45 nsew signal output
rlabel metal2 s 20160 100 20216 400 6 io_oeb[16]
port 46 nsew signal output
rlabel metal2 s 6720 100 6776 400 6 io_oeb[17]
port 47 nsew signal output
rlabel metal2 s 3360 69600 3416 69900 6 io_oeb[18]
port 48 nsew signal output
rlabel metal2 s 24864 69600 24920 69900 6 io_oeb[19]
port 49 nsew signal output
rlabel metal2 s 18816 69600 18872 69900 6 io_oeb[1]
port 50 nsew signal output
rlabel metal2 s 40320 69600 40376 69900 6 io_oeb[20]
port 51 nsew signal output
rlabel metal2 s 59808 100 59864 400 6 io_oeb[21]
port 52 nsew signal output
rlabel metal3 s 69600 18144 69900 18200 6 io_oeb[22]
port 53 nsew signal output
rlabel metal2 s 67872 69600 67928 69900 6 io_oeb[23]
port 54 nsew signal output
rlabel metal3 s 100 20160 400 20216 6 io_oeb[24]
port 55 nsew signal output
rlabel metal3 s 100 10080 400 10136 6 io_oeb[25]
port 56 nsew signal output
rlabel metal3 s 100 63840 400 63896 6 io_oeb[26]
port 57 nsew signal output
rlabel metal2 s 58464 100 58520 400 6 io_oeb[27]
port 58 nsew signal output
rlabel metal2 s 1344 69600 1400 69900 6 io_oeb[28]
port 59 nsew signal output
rlabel metal3 s 69600 35616 69900 35672 6 io_oeb[29]
port 60 nsew signal output
rlabel metal3 s 69600 26880 69900 26936 6 io_oeb[2]
port 61 nsew signal output
rlabel metal2 s 65856 100 65912 400 6 io_oeb[30]
port 62 nsew signal output
rlabel metal3 s 100 21504 400 21560 6 io_oeb[31]
port 63 nsew signal output
rlabel metal2 s 61152 69600 61208 69900 6 io_oeb[32]
port 64 nsew signal output
rlabel metal3 s 69600 11424 69900 11480 6 io_oeb[33]
port 65 nsew signal output
rlabel metal3 s 100 57120 400 57176 6 io_oeb[34]
port 66 nsew signal output
rlabel metal3 s 69600 63168 69900 63224 6 io_oeb[35]
port 67 nsew signal output
rlabel metal2 s 38976 69600 39032 69900 6 io_oeb[36]
port 68 nsew signal output
rlabel metal3 s 69600 28224 69900 28280 6 io_oeb[37]
port 69 nsew signal output
rlabel metal3 s 100 52416 400 52472 6 io_oeb[3]
port 70 nsew signal output
rlabel metal3 s 100 9408 400 9464 6 io_oeb[4]
port 71 nsew signal output
rlabel metal2 s 51072 69600 51128 69900 6 io_oeb[5]
port 72 nsew signal output
rlabel metal3 s 100 55104 400 55160 6 io_oeb[6]
port 73 nsew signal output
rlabel metal2 s 33600 69600 33656 69900 6 io_oeb[7]
port 74 nsew signal output
rlabel metal3 s 100 34944 400 35000 6 io_oeb[8]
port 75 nsew signal output
rlabel metal3 s 69600 67872 69900 67928 6 io_oeb[9]
port 76 nsew signal output
rlabel metal2 s 11424 69600 11480 69900 6 io_out[0]
port 77 nsew signal output
rlabel metal2 s 21504 69600 21560 69900 6 io_out[10]
port 78 nsew signal output
rlabel metal2 s 45024 100 45080 400 6 io_out[11]
port 79 nsew signal output
rlabel metal2 s 68544 69600 68600 69900 6 io_out[12]
port 80 nsew signal output
rlabel metal3 s 100 69888 400 69944 6 io_out[13]
port 81 nsew signal output
rlabel metal3 s 100 51744 400 51800 6 io_out[14]
port 82 nsew signal output
rlabel metal2 s 28224 100 28280 400 6 io_out[15]
port 83 nsew signal output
rlabel metal3 s 69600 58464 69900 58520 6 io_out[16]
port 84 nsew signal output
rlabel metal2 s 8064 100 8120 400 6 io_out[17]
port 85 nsew signal output
rlabel metal2 s 65184 100 65240 400 6 io_out[18]
port 86 nsew signal output
rlabel metal2 s 15456 69600 15512 69900 6 io_out[19]
port 87 nsew signal output
rlabel metal2 s 4704 100 4760 400 6 io_out[1]
port 88 nsew signal output
rlabel metal3 s 69600 6720 69900 6776 6 io_out[20]
port 89 nsew signal output
rlabel metal3 s 100 46368 400 46424 6 io_out[21]
port 90 nsew signal output
rlabel metal3 s 69600 15456 69900 15512 6 io_out[22]
port 91 nsew signal output
rlabel metal3 s 100 26208 400 26264 6 io_out[23]
port 92 nsew signal output
rlabel metal2 s 61152 100 61208 400 6 io_out[24]
port 93 nsew signal output
rlabel metal3 s 69600 2016 69900 2072 6 io_out[25]
port 94 nsew signal output
rlabel metal2 s 29568 100 29624 400 6 io_out[26]
port 95 nsew signal output
rlabel metal2 s 23520 100 23576 400 6 io_out[27]
port 96 nsew signal output
rlabel metal2 s 49056 69600 49112 69900 6 io_out[28]
port 97 nsew signal output
rlabel metal2 s 47712 100 47768 400 6 io_out[29]
port 98 nsew signal output
rlabel metal3 s 69600 24864 69900 24920 6 io_out[2]
port 99 nsew signal output
rlabel metal2 s 63840 69600 63896 69900 6 io_out[30]
port 100 nsew signal output
rlabel metal2 s 24864 100 24920 400 6 io_out[31]
port 101 nsew signal output
rlabel metal2 s 43680 69600 43736 69900 6 io_out[32]
port 102 nsew signal output
rlabel metal3 s 100 25536 400 25592 6 io_out[33]
port 103 nsew signal output
rlabel metal2 s 46368 100 46424 400 6 io_out[34]
port 104 nsew signal output
rlabel metal2 s 41664 100 41720 400 6 io_out[35]
port 105 nsew signal output
rlabel metal2 s 16800 100 16856 400 6 io_out[36]
port 106 nsew signal output
rlabel metal3 s 100 3360 400 3416 6 io_out[37]
port 107 nsew signal output
rlabel metal2 s 32256 69600 32312 69900 6 io_out[3]
port 108 nsew signal output
rlabel metal2 s 32256 100 32312 400 6 io_out[4]
port 109 nsew signal output
rlabel metal2 s 29568 69600 29624 69900 6 io_out[5]
port 110 nsew signal output
rlabel metal3 s 100 12768 400 12824 6 io_out[6]
port 111 nsew signal output
rlabel metal3 s 100 39648 400 39704 6 io_out[7]
port 112 nsew signal output
rlabel metal2 s 51072 100 51128 400 6 io_out[8]
port 113 nsew signal output
rlabel metal2 s 18144 100 18200 400 6 io_out[9]
port 114 nsew signal output
rlabel metal3 s 100 35616 400 35672 6 la_data_in[0]
port 115 nsew signal input
rlabel metal3 s 69600 65184 69900 65240 6 la_data_in[10]
port 116 nsew signal input
rlabel metal3 s 69600 30912 69900 30968 6 la_data_in[11]
port 117 nsew signal input
rlabel metal2 s 21504 100 21560 400 6 la_data_in[12]
port 118 nsew signal input
rlabel metal2 s 28224 69600 28280 69900 6 la_data_in[13]
port 119 nsew signal input
rlabel metal3 s 100 61152 400 61208 6 la_data_in[14]
port 120 nsew signal input
rlabel metal3 s 69600 50400 69900 50456 6 la_data_in[15]
port 121 nsew signal input
rlabel metal2 s 6720 69600 6776 69900 6 la_data_in[16]
port 122 nsew signal input
rlabel metal3 s 69600 10752 69900 10808 6 la_data_in[17]
port 123 nsew signal input
rlabel metal2 s 34944 69600 35000 69900 6 la_data_in[18]
port 124 nsew signal input
rlabel metal3 s 100 10752 400 10808 6 la_data_in[19]
port 125 nsew signal input
rlabel metal2 s 16128 69600 16184 69900 6 la_data_in[1]
port 126 nsew signal input
rlabel metal3 s 69600 14784 69900 14840 6 la_data_in[20]
port 127 nsew signal input
rlabel metal3 s 100 53088 400 53144 6 la_data_in[21]
port 128 nsew signal input
rlabel metal3 s 100 30912 400 30968 6 la_data_in[22]
port 129 nsew signal input
rlabel metal3 s 69600 52416 69900 52472 6 la_data_in[23]
port 130 nsew signal input
rlabel metal2 s 35616 69600 35672 69900 6 la_data_in[24]
port 131 nsew signal input
rlabel metal2 s 14784 69600 14840 69900 6 la_data_in[25]
port 132 nsew signal input
rlabel metal2 s 43008 69600 43064 69900 6 la_data_in[26]
port 133 nsew signal input
rlabel metal3 s 100 63168 400 63224 6 la_data_in[27]
port 134 nsew signal input
rlabel metal3 s 100 65856 400 65912 6 la_data_in[28]
port 135 nsew signal input
rlabel metal3 s 69600 17472 69900 17528 6 la_data_in[29]
port 136 nsew signal input
rlabel metal2 s 30912 69600 30968 69900 6 la_data_in[2]
port 137 nsew signal input
rlabel metal3 s 100 5376 400 5432 6 la_data_in[30]
port 138 nsew signal input
rlabel metal2 s 59136 69600 59192 69900 6 la_data_in[31]
port 139 nsew signal input
rlabel metal3 s 100 28224 400 28280 6 la_data_in[32]
port 140 nsew signal input
rlabel metal3 s 100 47040 400 47096 6 la_data_in[33]
port 141 nsew signal input
rlabel metal2 s 5376 69600 5432 69900 6 la_data_in[34]
port 142 nsew signal input
rlabel metal3 s 100 61824 400 61880 6 la_data_in[35]
port 143 nsew signal input
rlabel metal2 s 49728 100 49784 400 6 la_data_in[36]
port 144 nsew signal input
rlabel metal3 s 100 68544 400 68600 6 la_data_in[37]
port 145 nsew signal input
rlabel metal2 s 31584 100 31640 400 6 la_data_in[38]
port 146 nsew signal input
rlabel metal2 s 38304 69600 38360 69900 6 la_data_in[39]
port 147 nsew signal input
rlabel metal3 s 69600 38304 69900 38360 6 la_data_in[3]
port 148 nsew signal input
rlabel metal2 s 24192 100 24248 400 6 la_data_in[40]
port 149 nsew signal input
rlabel metal2 s 33600 100 33656 400 6 la_data_in[41]
port 150 nsew signal input
rlabel metal3 s 100 23520 400 23576 6 la_data_in[42]
port 151 nsew signal input
rlabel metal2 s 65856 69600 65912 69900 6 la_data_in[43]
port 152 nsew signal input
rlabel metal3 s 69600 672 69900 728 6 la_data_in[44]
port 153 nsew signal input
rlabel metal2 s 22848 100 22904 400 6 la_data_in[45]
port 154 nsew signal input
rlabel metal3 s 69600 51072 69900 51128 6 la_data_in[46]
port 155 nsew signal input
rlabel metal2 s 43680 100 43736 400 6 la_data_in[47]
port 156 nsew signal input
rlabel metal2 s 32928 69600 32984 69900 6 la_data_in[48]
port 157 nsew signal input
rlabel metal2 s 26880 69600 26936 69900 6 la_data_in[49]
port 158 nsew signal input
rlabel metal2 s 6048 69600 6104 69900 6 la_data_in[4]
port 159 nsew signal input
rlabel metal2 s 27552 69600 27608 69900 6 la_data_in[50]
port 160 nsew signal input
rlabel metal2 s 32928 100 32984 400 6 la_data_in[51]
port 161 nsew signal input
rlabel metal3 s 69600 23520 69900 23576 6 la_data_in[52]
port 162 nsew signal input
rlabel metal2 s 54432 69600 54488 69900 6 la_data_in[53]
port 163 nsew signal input
rlabel metal2 s 49728 69600 49784 69900 6 la_data_in[54]
port 164 nsew signal input
rlabel metal3 s 100 18816 400 18872 6 la_data_in[55]
port 165 nsew signal input
rlabel metal3 s 100 20832 400 20888 6 la_data_in[56]
port 166 nsew signal input
rlabel metal2 s 2016 69600 2072 69900 6 la_data_in[57]
port 167 nsew signal input
rlabel metal2 s 25536 100 25592 400 6 la_data_in[58]
port 168 nsew signal input
rlabel metal3 s 69600 63840 69900 63896 6 la_data_in[59]
port 169 nsew signal input
rlabel metal2 s 12096 100 12152 400 6 la_data_in[5]
port 170 nsew signal input
rlabel metal3 s 69600 46368 69900 46424 6 la_data_in[60]
port 171 nsew signal input
rlabel metal3 s 100 2016 400 2072 6 la_data_in[61]
port 172 nsew signal input
rlabel metal2 s 40992 100 41048 400 6 la_data_in[62]
port 173 nsew signal input
rlabel metal2 s 18144 69600 18200 69900 6 la_data_in[63]
port 174 nsew signal input
rlabel metal2 s 14112 100 14168 400 6 la_data_in[6]
port 175 nsew signal input
rlabel metal3 s 69600 25536 69900 25592 6 la_data_in[7]
port 176 nsew signal input
rlabel metal3 s 100 1344 400 1400 6 la_data_in[8]
port 177 nsew signal input
rlabel metal2 s 63168 69600 63224 69900 6 la_data_in[9]
port 178 nsew signal input
rlabel metal2 s 60480 69600 60536 69900 6 la_data_out[0]
port 179 nsew signal output
rlabel metal3 s 69600 37632 69900 37688 6 la_data_out[10]
port 180 nsew signal output
rlabel metal3 s 100 2688 400 2744 6 la_data_out[11]
port 181 nsew signal output
rlabel metal3 s 100 50400 400 50456 6 la_data_out[12]
port 182 nsew signal output
rlabel metal2 s 26208 100 26264 400 6 la_data_out[13]
port 183 nsew signal output
rlabel metal3 s 69600 28896 69900 28952 6 la_data_out[14]
port 184 nsew signal output
rlabel metal3 s 100 59808 400 59864 6 la_data_out[15]
port 185 nsew signal output
rlabel metal3 s 69600 38976 69900 39032 6 la_data_out[16]
port 186 nsew signal output
rlabel metal2 s 34272 69600 34328 69900 6 la_data_out[17]
port 187 nsew signal output
rlabel metal3 s 69600 57792 69900 57848 6 la_data_out[18]
port 188 nsew signal output
rlabel metal2 s 36960 100 37016 400 6 la_data_out[19]
port 189 nsew signal output
rlabel metal3 s 69600 32928 69900 32984 6 la_data_out[1]
port 190 nsew signal output
rlabel metal3 s 69600 10080 69900 10136 6 la_data_out[20]
port 191 nsew signal output
rlabel metal3 s 100 69216 400 69272 6 la_data_out[21]
port 192 nsew signal output
rlabel metal3 s 69600 43680 69900 43736 6 la_data_out[22]
port 193 nsew signal output
rlabel metal2 s 20832 100 20888 400 6 la_data_out[23]
port 194 nsew signal output
rlabel metal3 s 100 31584 400 31640 6 la_data_out[24]
port 195 nsew signal output
rlabel metal2 s 37632 100 37688 400 6 la_data_out[25]
port 196 nsew signal output
rlabel metal3 s 100 67872 400 67928 6 la_data_out[26]
port 197 nsew signal output
rlabel metal2 s 42336 69600 42392 69900 6 la_data_out[27]
port 198 nsew signal output
rlabel metal3 s 69600 55776 69900 55832 6 la_data_out[28]
port 199 nsew signal output
rlabel metal2 s 30240 100 30296 400 6 la_data_out[29]
port 200 nsew signal output
rlabel metal3 s 100 16128 400 16184 6 la_data_out[2]
port 201 nsew signal output
rlabel metal3 s 69600 32256 69900 32312 6 la_data_out[30]
port 202 nsew signal output
rlabel metal3 s 69600 3360 69900 3416 6 la_data_out[31]
port 203 nsew signal output
rlabel metal2 s 40992 69600 41048 69900 6 la_data_out[32]
port 204 nsew signal output
rlabel metal3 s 69600 12768 69900 12824 6 la_data_out[33]
port 205 nsew signal output
rlabel metal2 s 34272 100 34328 400 6 la_data_out[34]
port 206 nsew signal output
rlabel metal2 s 37632 69600 37688 69900 6 la_data_out[35]
port 207 nsew signal output
rlabel metal3 s 69600 56448 69900 56504 6 la_data_out[36]
port 208 nsew signal output
rlabel metal3 s 69600 27552 69900 27608 6 la_data_out[37]
port 209 nsew signal output
rlabel metal3 s 69600 1344 69900 1400 6 la_data_out[38]
port 210 nsew signal output
rlabel metal3 s 69600 9408 69900 9464 6 la_data_out[39]
port 211 nsew signal output
rlabel metal3 s 100 11424 400 11480 6 la_data_out[3]
port 212 nsew signal output
rlabel metal2 s 67872 100 67928 400 6 la_data_out[40]
port 213 nsew signal output
rlabel metal3 s 69600 21504 69900 21560 6 la_data_out[41]
port 214 nsew signal output
rlabel metal3 s 69600 59136 69900 59192 6 la_data_out[42]
port 215 nsew signal output
rlabel metal2 s 4032 100 4088 400 6 la_data_out[43]
port 216 nsew signal output
rlabel metal2 s 28896 100 28952 400 6 la_data_out[44]
port 217 nsew signal output
rlabel metal2 s 10752 69600 10808 69900 6 la_data_out[45]
port 218 nsew signal output
rlabel metal2 s 10080 69600 10136 69900 6 la_data_out[46]
port 219 nsew signal output
rlabel metal3 s 100 49728 400 49784 6 la_data_out[47]
port 220 nsew signal output
rlabel metal2 s 16128 100 16184 400 6 la_data_out[48]
port 221 nsew signal output
rlabel metal2 s 63168 100 63224 400 6 la_data_out[49]
port 222 nsew signal output
rlabel metal2 s 39648 69600 39704 69900 6 la_data_out[4]
port 223 nsew signal output
rlabel metal2 s 24192 69600 24248 69900 6 la_data_out[50]
port 224 nsew signal output
rlabel metal3 s 100 67200 400 67256 6 la_data_out[51]
port 225 nsew signal output
rlabel metal3 s 69600 4704 69900 4760 6 la_data_out[52]
port 226 nsew signal output
rlabel metal3 s 100 66528 400 66584 6 la_data_out[53]
port 227 nsew signal output
rlabel metal3 s 69600 47712 69900 47768 6 la_data_out[54]
port 228 nsew signal output
rlabel metal2 s 26208 69600 26264 69900 6 la_data_out[55]
port 229 nsew signal output
rlabel metal3 s 69600 16800 69900 16856 6 la_data_out[56]
port 230 nsew signal output
rlabel metal2 s 53088 69600 53144 69900 6 la_data_out[57]
port 231 nsew signal output
rlabel metal3 s 69600 48384 69900 48440 6 la_data_out[58]
port 232 nsew signal output
rlabel metal3 s 100 26880 400 26936 6 la_data_out[59]
port 233 nsew signal output
rlabel metal3 s 69600 41664 69900 41720 6 la_data_out[5]
port 234 nsew signal output
rlabel metal2 s 56448 69600 56504 69900 6 la_data_out[60]
port 235 nsew signal output
rlabel metal2 s 18816 100 18872 400 6 la_data_out[61]
port 236 nsew signal output
rlabel metal2 s 60480 100 60536 400 6 la_data_out[62]
port 237 nsew signal output
rlabel metal3 s 69600 5376 69900 5432 6 la_data_out[63]
port 238 nsew signal output
rlabel metal3 s 69600 20160 69900 20216 6 la_data_out[6]
port 239 nsew signal output
rlabel metal2 s 67200 69600 67256 69900 6 la_data_out[7]
port 240 nsew signal output
rlabel metal3 s 100 4032 400 4088 6 la_data_out[8]
port 241 nsew signal output
rlabel metal3 s 69600 33600 69900 33656 6 la_data_out[9]
port 242 nsew signal output
rlabel metal3 s 69600 26208 69900 26264 6 la_oenb[0]
port 243 nsew signal input
rlabel metal3 s 69600 49728 69900 49784 6 la_oenb[10]
port 244 nsew signal input
rlabel metal3 s 69600 39648 69900 39704 6 la_oenb[11]
port 245 nsew signal input
rlabel metal2 s 672 69600 728 69900 6 la_oenb[12]
port 246 nsew signal input
rlabel metal3 s 100 55776 400 55832 6 la_oenb[13]
port 247 nsew signal input
rlabel metal2 s 51744 100 51800 400 6 la_oenb[14]
port 248 nsew signal input
rlabel metal2 s 61824 100 61880 400 6 la_oenb[15]
port 249 nsew signal input
rlabel metal2 s 10080 100 10136 400 6 la_oenb[16]
port 250 nsew signal input
rlabel metal3 s 100 8736 400 8792 6 la_oenb[17]
port 251 nsew signal input
rlabel metal2 s 4704 69600 4760 69900 6 la_oenb[18]
port 252 nsew signal input
rlabel metal3 s 69600 6048 69900 6104 6 la_oenb[19]
port 253 nsew signal input
rlabel metal2 s 13440 69600 13496 69900 6 la_oenb[1]
port 254 nsew signal input
rlabel metal3 s 100 40992 400 41048 6 la_oenb[20]
port 255 nsew signal input
rlabel metal2 s 28896 69600 28952 69900 6 la_oenb[21]
port 256 nsew signal input
rlabel metal2 s 51744 69600 51800 69900 6 la_oenb[22]
port 257 nsew signal input
rlabel metal2 s 19488 100 19544 400 6 la_oenb[23]
port 258 nsew signal input
rlabel metal3 s 69600 43008 69900 43064 6 la_oenb[24]
port 259 nsew signal input
rlabel metal2 s 62496 100 62552 400 6 la_oenb[25]
port 260 nsew signal input
rlabel metal2 s 14112 69600 14168 69900 6 la_oenb[26]
port 261 nsew signal input
rlabel metal2 s 12768 100 12824 400 6 la_oenb[27]
port 262 nsew signal input
rlabel metal3 s 100 43008 400 43064 6 la_oenb[28]
port 263 nsew signal input
rlabel metal3 s 69600 66528 69900 66584 6 la_oenb[29]
port 264 nsew signal input
rlabel metal2 s 69216 69600 69272 69900 6 la_oenb[2]
port 265 nsew signal input
rlabel metal3 s 69600 59808 69900 59864 6 la_oenb[30]
port 266 nsew signal input
rlabel metal2 s 30240 69600 30296 69900 6 la_oenb[31]
port 267 nsew signal input
rlabel metal3 s 69600 57120 69900 57176 6 la_oenb[32]
port 268 nsew signal input
rlabel metal2 s 35616 100 35672 400 6 la_oenb[33]
port 269 nsew signal input
rlabel metal2 s 12096 69600 12152 69900 6 la_oenb[34]
port 270 nsew signal input
rlabel metal2 s 2016 100 2072 400 6 la_oenb[35]
port 271 nsew signal input
rlabel metal2 s 672 100 728 400 6 la_oenb[36]
port 272 nsew signal input
rlabel metal2 s 9408 69600 9464 69900 6 la_oenb[37]
port 273 nsew signal input
rlabel metal2 s 36288 100 36344 400 6 la_oenb[38]
port 274 nsew signal input
rlabel metal3 s 100 30240 400 30296 6 la_oenb[39]
port 275 nsew signal input
rlabel metal3 s 100 38304 400 38360 6 la_oenb[3]
port 276 nsew signal input
rlabel metal3 s 69600 8736 69900 8792 6 la_oenb[40]
port 277 nsew signal input
rlabel metal2 s 25536 69600 25592 69900 6 la_oenb[41]
port 278 nsew signal input
rlabel metal3 s 100 44352 400 44408 6 la_oenb[42]
port 279 nsew signal input
rlabel metal2 s 13440 100 13496 400 6 la_oenb[43]
port 280 nsew signal input
rlabel metal2 s 30912 100 30968 400 6 la_oenb[44]
port 281 nsew signal input
rlabel metal2 s 57792 69600 57848 69900 6 la_oenb[45]
port 282 nsew signal input
rlabel metal2 s 55776 100 55832 400 6 la_oenb[46]
port 283 nsew signal input
rlabel metal3 s 100 8064 400 8120 6 la_oenb[47]
port 284 nsew signal input
rlabel metal3 s 100 51072 400 51128 6 la_oenb[48]
port 285 nsew signal input
rlabel metal3 s 100 672 400 728 6 la_oenb[49]
port 286 nsew signal input
rlabel metal3 s 100 65184 400 65240 6 la_oenb[4]
port 287 nsew signal input
rlabel metal2 s 53760 100 53816 400 6 la_oenb[50]
port 288 nsew signal input
rlabel metal2 s 22848 69600 22904 69900 6 la_oenb[51]
port 289 nsew signal input
rlabel metal2 s 69216 100 69272 400 6 la_oenb[52]
port 290 nsew signal input
rlabel metal3 s 69600 44352 69900 44408 6 la_oenb[53]
port 291 nsew signal input
rlabel metal3 s 100 37632 400 37688 6 la_oenb[54]
port 292 nsew signal input
rlabel metal3 s 69600 36288 69900 36344 6 la_oenb[55]
port 293 nsew signal input
rlabel metal2 s 53088 100 53144 400 6 la_oenb[56]
port 294 nsew signal input
rlabel metal2 s 61824 69600 61880 69900 6 la_oenb[57]
port 295 nsew signal input
rlabel metal3 s 69600 7392 69900 7448 6 la_oenb[58]
port 296 nsew signal input
rlabel metal2 s 41664 69600 41720 69900 6 la_oenb[59]
port 297 nsew signal input
rlabel metal2 s 64512 100 64568 400 6 la_oenb[5]
port 298 nsew signal input
rlabel metal3 s 100 34272 400 34328 6 la_oenb[60]
port 299 nsew signal input
rlabel metal2 s 8736 100 8792 400 6 la_oenb[61]
port 300 nsew signal input
rlabel metal3 s 69600 34944 69900 35000 6 la_oenb[62]
port 301 nsew signal input
rlabel metal3 s 100 16800 400 16856 6 la_oenb[63]
port 302 nsew signal input
rlabel metal3 s 69600 45696 69900 45752 6 la_oenb[6]
port 303 nsew signal input
rlabel metal2 s 17472 100 17528 400 6 la_oenb[7]
port 304 nsew signal input
rlabel metal2 s 66528 100 66584 400 6 la_oenb[8]
port 305 nsew signal input
rlabel metal2 s 20160 69600 20216 69900 6 la_oenb[9]
port 306 nsew signal input
rlabel metal2 s 59808 69600 59864 69900 6 user_clock2
port 307 nsew signal input
rlabel metal3 s 69600 53760 69900 53816 6 user_irq[0]
port 308 nsew signal output
rlabel metal2 s 17472 69600 17528 69900 6 user_irq[1]
port 309 nsew signal output
rlabel metal3 s 100 45024 400 45080 6 user_irq[2]
port 310 nsew signal output
rlabel metal4 s 2224 1538 2384 68238 6 vdd
port 311 nsew power bidirectional
rlabel metal4 s 17584 1538 17744 68238 6 vdd
port 311 nsew power bidirectional
rlabel metal4 s 32944 1538 33104 68238 6 vdd
port 311 nsew power bidirectional
rlabel metal4 s 48304 1538 48464 68238 6 vdd
port 311 nsew power bidirectional
rlabel metal4 s 63664 1538 63824 68238 6 vdd
port 311 nsew power bidirectional
rlabel metal4 s 9904 1538 10064 68238 6 vss
port 312 nsew ground bidirectional
rlabel metal4 s 25264 1538 25424 68238 6 vss
port 312 nsew ground bidirectional
rlabel metal4 s 40624 1538 40784 68238 6 vss
port 312 nsew ground bidirectional
rlabel metal4 s 55984 1538 56144 68238 6 vss
port 312 nsew ground bidirectional
rlabel metal3 s 69600 12096 69900 12152 6 wb_clk_i
port 313 nsew signal input
rlabel metal2 s 12768 69600 12824 69900 6 wb_rst_i
port 314 nsew signal input
rlabel metal3 s 69600 24192 69900 24248 6 wbs_ack_o
port 315 nsew signal output
rlabel metal2 s 46368 69600 46424 69900 6 wbs_adr_i[0]
port 316 nsew signal input
rlabel metal2 s 31584 69600 31640 69900 6 wbs_adr_i[10]
port 317 nsew signal input
rlabel metal3 s 100 40320 400 40376 6 wbs_adr_i[11]
port 318 nsew signal input
rlabel metal2 s 6048 100 6104 400 6 wbs_adr_i[12]
port 319 nsew signal input
rlabel metal2 s 38976 100 39032 400 6 wbs_adr_i[13]
port 320 nsew signal input
rlabel metal3 s 100 6720 400 6776 6 wbs_adr_i[14]
port 321 nsew signal input
rlabel metal3 s 69600 47040 69900 47096 6 wbs_adr_i[15]
port 322 nsew signal input
rlabel metal2 s 44352 100 44408 400 6 wbs_adr_i[16]
port 323 nsew signal input
rlabel metal3 s 100 38976 400 39032 6 wbs_adr_i[17]
port 324 nsew signal input
rlabel metal3 s 69600 22176 69900 22232 6 wbs_adr_i[18]
port 325 nsew signal input
rlabel metal2 s 67200 100 67256 400 6 wbs_adr_i[19]
port 326 nsew signal input
rlabel metal3 s 100 4704 400 4760 6 wbs_adr_i[1]
port 327 nsew signal input
rlabel metal2 s 65184 69600 65240 69900 6 wbs_adr_i[20]
port 328 nsew signal input
rlabel metal2 s 39648 100 39704 400 6 wbs_adr_i[21]
port 329 nsew signal input
rlabel metal2 s 56448 100 56504 400 6 wbs_adr_i[22]
port 330 nsew signal input
rlabel metal3 s 69600 16128 69900 16184 6 wbs_adr_i[23]
port 331 nsew signal input
rlabel metal2 s 8064 69600 8120 69900 6 wbs_adr_i[24]
port 332 nsew signal input
rlabel metal3 s 100 12096 400 12152 6 wbs_adr_i[25]
port 333 nsew signal input
rlabel metal2 s 7392 100 7448 400 6 wbs_adr_i[26]
port 334 nsew signal input
rlabel metal2 s 23520 69600 23576 69900 6 wbs_adr_i[27]
port 335 nsew signal input
rlabel metal3 s 69600 40992 69900 41048 6 wbs_adr_i[28]
port 336 nsew signal input
rlabel metal3 s 69600 67200 69900 67256 6 wbs_adr_i[29]
port 337 nsew signal input
rlabel metal2 s 27552 100 27608 400 6 wbs_adr_i[2]
port 338 nsew signal input
rlabel metal3 s 100 27552 400 27608 6 wbs_adr_i[30]
port 339 nsew signal input
rlabel metal3 s 69600 29568 69900 29624 6 wbs_adr_i[31]
port 340 nsew signal input
rlabel metal2 s 54432 100 54488 400 6 wbs_adr_i[3]
port 341 nsew signal input
rlabel metal2 s 53760 69600 53816 69900 6 wbs_adr_i[4]
port 342 nsew signal input
rlabel metal2 s 52416 100 52472 400 6 wbs_adr_i[5]
port 343 nsew signal input
rlabel metal3 s 100 17472 400 17528 6 wbs_adr_i[6]
port 344 nsew signal input
rlabel metal2 s 3360 100 3416 400 6 wbs_adr_i[7]
port 345 nsew signal input
rlabel metal3 s 69600 0 69900 56 6 wbs_adr_i[8]
port 346 nsew signal input
rlabel metal3 s 69600 18816 69900 18872 6 wbs_adr_i[9]
port 347 nsew signal input
rlabel metal2 s 22176 69600 22232 69900 6 wbs_cyc_i
port 348 nsew signal input
rlabel metal3 s 69600 61152 69900 61208 6 wbs_dat_i[0]
port 349 nsew signal input
rlabel metal3 s 100 53760 400 53816 6 wbs_dat_i[10]
port 350 nsew signal input
rlabel metal3 s 100 59136 400 59192 6 wbs_dat_i[11]
port 351 nsew signal input
rlabel metal3 s 100 56448 400 56504 6 wbs_dat_i[12]
port 352 nsew signal input
rlabel metal2 s 2688 100 2744 400 6 wbs_dat_i[13]
port 353 nsew signal input
rlabel metal3 s 100 14784 400 14840 6 wbs_dat_i[14]
port 354 nsew signal input
rlabel metal3 s 69600 36960 69900 37016 6 wbs_dat_i[15]
port 355 nsew signal input
rlabel metal2 s 40320 100 40376 400 6 wbs_dat_i[16]
port 356 nsew signal input
rlabel metal2 s 47712 69600 47768 69900 6 wbs_dat_i[17]
port 357 nsew signal input
rlabel metal2 s 64512 69600 64568 69900 6 wbs_dat_i[18]
port 358 nsew signal input
rlabel metal2 s 4032 69600 4088 69900 6 wbs_dat_i[19]
port 359 nsew signal input
rlabel metal2 s 10752 100 10808 400 6 wbs_dat_i[1]
port 360 nsew signal input
rlabel metal3 s 100 32928 400 32984 6 wbs_dat_i[20]
port 361 nsew signal input
rlabel metal2 s 66528 69600 66584 69900 6 wbs_dat_i[21]
port 362 nsew signal input
rlabel metal3 s 100 41664 400 41720 6 wbs_dat_i[22]
port 363 nsew signal input
rlabel metal3 s 69600 55104 69900 55160 6 wbs_dat_i[23]
port 364 nsew signal input
rlabel metal3 s 69600 22848 69900 22904 6 wbs_dat_i[24]
port 365 nsew signal input
rlabel metal2 s 48384 100 48440 400 6 wbs_dat_i[25]
port 366 nsew signal input
rlabel metal2 s 58464 69600 58520 69900 6 wbs_dat_i[26]
port 367 nsew signal input
rlabel metal2 s 16800 69600 16856 69900 6 wbs_dat_i[27]
port 368 nsew signal input
rlabel metal2 s 22176 100 22232 400 6 wbs_dat_i[28]
port 369 nsew signal input
rlabel metal3 s 69600 42336 69900 42392 6 wbs_dat_i[29]
port 370 nsew signal input
rlabel metal2 s 57120 100 57176 400 6 wbs_dat_i[2]
port 371 nsew signal input
rlabel metal3 s 69600 20832 69900 20888 6 wbs_dat_i[30]
port 372 nsew signal input
rlabel metal3 s 100 36960 400 37016 6 wbs_dat_i[31]
port 373 nsew signal input
rlabel metal3 s 69600 2688 69900 2744 6 wbs_dat_i[3]
port 374 nsew signal input
rlabel metal2 s 11424 100 11480 400 6 wbs_dat_i[4]
port 375 nsew signal input
rlabel metal2 s 34944 100 35000 400 6 wbs_dat_i[5]
port 376 nsew signal input
rlabel metal3 s 69600 30240 69900 30296 6 wbs_dat_i[6]
port 377 nsew signal input
rlabel metal2 s 55104 69600 55160 69900 6 wbs_dat_i[7]
port 378 nsew signal input
rlabel metal3 s 69600 62496 69900 62552 6 wbs_dat_i[8]
port 379 nsew signal input
rlabel metal3 s 69600 4032 69900 4088 6 wbs_dat_i[9]
port 380 nsew signal input
rlabel metal3 s 100 14112 400 14168 6 wbs_dat_o[0]
port 381 nsew signal output
rlabel metal3 s 69600 40320 69900 40376 6 wbs_dat_o[10]
port 382 nsew signal output
rlabel metal2 s 1344 100 1400 400 6 wbs_dat_o[11]
port 383 nsew signal output
rlabel metal3 s 69600 64512 69900 64568 6 wbs_dat_o[12]
port 384 nsew signal output
rlabel metal2 s 52416 69600 52472 69900 6 wbs_dat_o[13]
port 385 nsew signal output
rlabel metal3 s 69600 8064 69900 8120 6 wbs_dat_o[14]
port 386 nsew signal output
rlabel metal2 s 50400 69600 50456 69900 6 wbs_dat_o[15]
port 387 nsew signal output
rlabel metal3 s 100 19488 400 19544 6 wbs_dat_o[16]
port 388 nsew signal output
rlabel metal3 s 100 22176 400 22232 6 wbs_dat_o[17]
port 389 nsew signal output
rlabel metal2 s 47040 100 47096 400 6 wbs_dat_o[18]
port 390 nsew signal output
rlabel metal2 s 0 100 56 400 6 wbs_dat_o[19]
port 391 nsew signal output
rlabel metal2 s 55104 100 55160 400 6 wbs_dat_o[1]
port 392 nsew signal output
rlabel metal3 s 100 33600 400 33656 6 wbs_dat_o[20]
port 393 nsew signal output
rlabel metal3 s 100 60480 400 60536 6 wbs_dat_o[21]
port 394 nsew signal output
rlabel metal2 s 19488 69600 19544 69900 6 wbs_dat_o[22]
port 395 nsew signal output
rlabel metal3 s 100 22848 400 22904 6 wbs_dat_o[23]
port 396 nsew signal output
rlabel metal2 s 14784 100 14840 400 6 wbs_dat_o[24]
port 397 nsew signal output
rlabel metal2 s 5376 100 5432 400 6 wbs_dat_o[25]
port 398 nsew signal output
rlabel metal2 s 36288 69600 36344 69900 6 wbs_dat_o[26]
port 399 nsew signal output
rlabel metal2 s 20832 69600 20888 69900 6 wbs_dat_o[27]
port 400 nsew signal output
rlabel metal2 s 38304 100 38360 400 6 wbs_dat_o[28]
port 401 nsew signal output
rlabel metal2 s 48384 69600 48440 69900 6 wbs_dat_o[29]
port 402 nsew signal output
rlabel metal3 s 69600 19488 69900 19544 6 wbs_dat_o[2]
port 403 nsew signal output
rlabel metal3 s 100 45696 400 45752 6 wbs_dat_o[30]
port 404 nsew signal output
rlabel metal3 s 69600 54432 69900 54488 6 wbs_dat_o[31]
port 405 nsew signal output
rlabel metal2 s 15456 100 15512 400 6 wbs_dat_o[3]
port 406 nsew signal output
rlabel metal2 s 26880 100 26936 400 6 wbs_dat_o[4]
port 407 nsew signal output
rlabel metal3 s 100 6048 400 6104 6 wbs_dat_o[5]
port 408 nsew signal output
rlabel metal3 s 69600 51744 69900 51800 6 wbs_dat_o[6]
port 409 nsew signal output
rlabel metal2 s 42336 100 42392 400 6 wbs_dat_o[7]
port 410 nsew signal output
rlabel metal2 s 45696 69600 45752 69900 6 wbs_dat_o[8]
port 411 nsew signal output
rlabel metal2 s 45024 69600 45080 69900 6 wbs_dat_o[9]
port 412 nsew signal output
rlabel metal3 s 100 64512 400 64568 6 wbs_sel_i[0]
port 413 nsew signal input
rlabel metal2 s 7392 69600 7448 69900 6 wbs_sel_i[1]
port 414 nsew signal input
rlabel metal2 s 50400 100 50456 400 6 wbs_sel_i[2]
port 415 nsew signal input
rlabel metal3 s 100 15456 400 15512 6 wbs_sel_i[3]
port 416 nsew signal input
rlabel metal3 s 100 57792 400 57848 6 wbs_stb_i
port 417 nsew signal input
rlabel metal3 s 69600 34272 69900 34328 6 wbs_we_i
port 418 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 70000 70000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 11816614
string GDS_FILE /home/runner/work/tiny_user_project_RISCV_with_CNN_coprocessor/tiny_user_project_RISCV_with_CNN_coprocessor/openlane/tiny_user_project/runs/22_12_02_17_21/results/signoff/tiny_user_project.magic.gds
string GDS_START 352256
<< end >>

